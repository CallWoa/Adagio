module Manager(
  input          clock,
  input          reset,
  input          io_mixPc, // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 135:14]
  input          io_uart_ctrl_tx_done, // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 135:14]
  input          io_uart_ctrl_rx_valid, // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 135:14]
  output         io_uart_ctrl_tx_en, // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 135:14]
  input          io_uart_rf_w_en, // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 135:14]
  input  [7:0]   io_uart_rf_r_addr, // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 135:14]
  input  [7:0]   io_uart_rf_w_addr, // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 135:14]
  output [63:0]  io_uart_rf_r_data, // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 135:14]
  input  [63:0]  io_uart_rf_w_data, // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 135:14]
  input          io_top_src_ready, // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 135:14]
  output         io_top_src_valid, // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 135:14]
  output [255:0] io_top_src_bits_tc0_ot0_tg0_matrix_a, // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 135:14]
  output [255:0] io_top_src_bits_tc0_ot0_tg0_matrix_b, // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 135:14]
  output [255:0] io_top_src_bits_tc0_ot0_tg0_matrix_c, // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 135:14]
  output [255:0] io_top_src_bits_tc0_ot0_tg4_matrix_a, // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 135:14]
  output [255:0] io_top_src_bits_tc0_ot0_tg4_matrix_b, // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 135:14]
  output [255:0] io_top_src_bits_tc0_ot0_tg4_matrix_c, // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 135:14]
  output [255:0] io_top_src_bits_tc0_ot1_tg0_matrix_a, // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 135:14]
  output [255:0] io_top_src_bits_tc0_ot1_tg0_matrix_b, // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 135:14]
  output [255:0] io_top_src_bits_tc0_ot1_tg0_matrix_c, // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 135:14]
  output [255:0] io_top_src_bits_tc0_ot1_tg4_matrix_a, // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 135:14]
  output [255:0] io_top_src_bits_tc0_ot1_tg4_matrix_b, // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 135:14]
  output [255:0] io_top_src_bits_tc0_ot1_tg4_matrix_c, // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 135:14]
  output [255:0] io_top_src_bits_tc1_ot0_tg0_matrix_a, // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 135:14]
  output [255:0] io_top_src_bits_tc1_ot0_tg0_matrix_b, // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 135:14]
  output [255:0] io_top_src_bits_tc1_ot0_tg0_matrix_c, // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 135:14]
  output [255:0] io_top_src_bits_tc1_ot0_tg4_matrix_a, // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 135:14]
  output [255:0] io_top_src_bits_tc1_ot0_tg4_matrix_b, // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 135:14]
  output [255:0] io_top_src_bits_tc1_ot0_tg4_matrix_c, // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 135:14]
  output [255:0] io_top_src_bits_tc1_ot1_tg0_matrix_a, // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 135:14]
  output [255:0] io_top_src_bits_tc1_ot1_tg0_matrix_b, // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 135:14]
  output [255:0] io_top_src_bits_tc1_ot1_tg0_matrix_c, // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 135:14]
  output [255:0] io_top_src_bits_tc1_ot1_tg4_matrix_a, // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 135:14]
  output [255:0] io_top_src_bits_tc1_ot1_tg4_matrix_b, // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 135:14]
  output [255:0] io_top_src_bits_tc1_ot1_tg4_matrix_c, // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 135:14]
  output         io_top_src_bits_ctrl_matBSel, // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 135:14]
  output         io_top_src_bits_ctrl_mixPcMode, // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 135:14]
  output         io_top_wb_ready, // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 135:14]
  input          io_top_wb_valid, // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 135:14]
  input  [255:0] io_top_wb_bits_tc0_octet0_threadgroup0_matrix_d_data, // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 135:14]
  input  [255:0] io_top_wb_bits_tc0_octet0_threadgroup4_matrix_d_data, // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 135:14]
  input  [255:0] io_top_wb_bits_tc0_octet1_threadgroup0_matrix_d_data, // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 135:14]
  input  [255:0] io_top_wb_bits_tc0_octet1_threadgroup4_matrix_d_data, // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 135:14]
  input  [255:0] io_top_wb_bits_tc1_octet0_threadgroup0_matrix_d_data, // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 135:14]
  input  [255:0] io_top_wb_bits_tc1_octet0_threadgroup4_matrix_d_data, // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 135:14]
  input  [255:0] io_top_wb_bits_tc1_octet1_threadgroup0_matrix_d_data, // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 135:14]
  input  [255:0] io_top_wb_bits_tc1_octet1_threadgroup4_matrix_d_data // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 135:14]
);
`ifdef RANDOMIZE_MEM_INIT
  reg [63:0] _RAND_0;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [255:0] _RAND_7;
  reg [255:0] _RAND_8;
  reg [255:0] _RAND_9;
  reg [255:0] _RAND_10;
  reg [255:0] _RAND_11;
  reg [255:0] _RAND_12;
  reg [255:0] _RAND_13;
  reg [255:0] _RAND_14;
  reg [255:0] _RAND_15;
  reg [255:0] _RAND_16;
  reg [255:0] _RAND_17;
  reg [255:0] _RAND_18;
  reg [255:0] _RAND_19;
  reg [255:0] _RAND_20;
  reg [255:0] _RAND_21;
  reg [255:0] _RAND_22;
  reg [255:0] _RAND_23;
  reg [255:0] _RAND_24;
  reg [255:0] _RAND_25;
  reg [255:0] _RAND_26;
  reg [255:0] _RAND_27;
  reg [255:0] _RAND_28;
  reg [255:0] _RAND_29;
  reg [255:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
`endif // RANDOMIZE_REG_INIT
  reg [63:0] rf [0:255]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_1_MPORT_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_1_MPORT_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_1_MPORT_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_0_MPORT_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_0_MPORT_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_0_MPORT_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_0_tile_v_3_MPORT_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_0_tile_v_3_MPORT_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_0_tile_v_3_MPORT_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_0_tile_v_2_MPORT_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_0_tile_v_2_MPORT_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_0_tile_v_2_MPORT_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_0_tile_v_1_MPORT_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_0_tile_v_1_MPORT_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_0_tile_v_1_MPORT_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_0_tile_v_0_MPORT_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_0_tile_v_0_MPORT_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_0_tile_v_0_MPORT_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_0_tile_v_3_MPORT_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_0_tile_v_3_MPORT_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_0_tile_v_3_MPORT_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_0_tile_v_2_MPORT_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_0_tile_v_2_MPORT_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_0_tile_v_2_MPORT_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_0_tile_v_1_MPORT_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_0_tile_v_1_MPORT_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_0_tile_v_1_MPORT_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_0_tile_v_0_MPORT_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_0_tile_v_0_MPORT_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_0_tile_v_0_MPORT_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_3_MPORT_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_3_MPORT_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_3_MPORT_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_2_MPORT_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_2_MPORT_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_2_MPORT_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_1_MPORT_1_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_1_MPORT_1_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_1_MPORT_1_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_0_MPORT_1_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_0_MPORT_1_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_0_MPORT_1_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_0_tile_v_3_MPORT_1_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_0_tile_v_3_MPORT_1_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_0_tile_v_3_MPORT_1_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_0_tile_v_2_MPORT_1_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_0_tile_v_2_MPORT_1_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_0_tile_v_2_MPORT_1_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_0_tile_v_1_MPORT_1_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_0_tile_v_1_MPORT_1_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_0_tile_v_1_MPORT_1_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_0_tile_v_0_MPORT_1_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_0_tile_v_0_MPORT_1_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_0_tile_v_0_MPORT_1_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_0_tile_v_3_MPORT_1_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_0_tile_v_3_MPORT_1_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_0_tile_v_3_MPORT_1_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_0_tile_v_2_MPORT_1_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_0_tile_v_2_MPORT_1_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_0_tile_v_2_MPORT_1_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_0_tile_v_1_MPORT_1_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_0_tile_v_1_MPORT_1_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_0_tile_v_1_MPORT_1_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_0_tile_v_0_MPORT_1_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_0_tile_v_0_MPORT_1_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_0_tile_v_0_MPORT_1_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_1_MPORT_2_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_1_MPORT_2_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_1_MPORT_2_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_0_MPORT_2_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_0_MPORT_2_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_0_MPORT_2_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_0_tile_v_3_MPORT_2_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_0_tile_v_3_MPORT_2_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_0_tile_v_3_MPORT_2_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_0_tile_v_2_MPORT_2_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_0_tile_v_2_MPORT_2_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_0_tile_v_2_MPORT_2_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_0_tile_v_1_MPORT_2_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_0_tile_v_1_MPORT_2_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_0_tile_v_1_MPORT_2_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_0_tile_v_0_MPORT_2_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_0_tile_v_0_MPORT_2_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_0_tile_v_0_MPORT_2_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_0_tile_v_3_MPORT_2_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_0_tile_v_3_MPORT_2_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_0_tile_v_3_MPORT_2_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_0_tile_v_2_MPORT_2_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_0_tile_v_2_MPORT_2_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_0_tile_v_2_MPORT_2_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_0_tile_v_1_MPORT_2_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_0_tile_v_1_MPORT_2_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_0_tile_v_1_MPORT_2_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_0_tile_v_0_MPORT_2_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_0_tile_v_0_MPORT_2_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_0_tile_v_0_MPORT_2_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_3_MPORT_1_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_3_MPORT_1_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_3_MPORT_1_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_2_MPORT_1_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_2_MPORT_1_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_2_MPORT_1_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_1_MPORT_3_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_1_MPORT_3_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_1_MPORT_3_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_0_MPORT_3_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_0_MPORT_3_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_0_MPORT_3_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_0_tile_v_3_MPORT_3_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_0_tile_v_3_MPORT_3_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_0_tile_v_3_MPORT_3_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_0_tile_v_2_MPORT_3_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_0_tile_v_2_MPORT_3_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_0_tile_v_2_MPORT_3_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_0_tile_v_1_MPORT_3_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_0_tile_v_1_MPORT_3_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_0_tile_v_1_MPORT_3_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_0_tile_v_0_MPORT_3_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_0_tile_v_0_MPORT_3_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_0_tile_v_0_MPORT_3_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_0_tile_v_3_MPORT_3_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_0_tile_v_3_MPORT_3_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_0_tile_v_3_MPORT_3_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_0_tile_v_2_MPORT_3_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_0_tile_v_2_MPORT_3_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_0_tile_v_2_MPORT_3_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_0_tile_v_1_MPORT_3_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_0_tile_v_1_MPORT_3_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_0_tile_v_1_MPORT_3_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_0_tile_v_0_MPORT_3_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_0_tile_v_0_MPORT_3_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_0_tile_v_0_MPORT_3_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_1_MPORT_4_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_1_MPORT_4_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_1_MPORT_4_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_0_MPORT_4_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_0_MPORT_4_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_0_MPORT_4_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_0_tile_v_3_MPORT_4_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_0_tile_v_3_MPORT_4_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_0_tile_v_3_MPORT_4_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_0_tile_v_2_MPORT_4_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_0_tile_v_2_MPORT_4_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_0_tile_v_2_MPORT_4_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_0_tile_v_1_MPORT_4_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_0_tile_v_1_MPORT_4_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_0_tile_v_1_MPORT_4_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_0_tile_v_0_MPORT_4_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_0_tile_v_0_MPORT_4_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_0_tile_v_0_MPORT_4_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_0_tile_v_3_MPORT_4_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_0_tile_v_3_MPORT_4_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_0_tile_v_3_MPORT_4_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_0_tile_v_2_MPORT_4_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_0_tile_v_2_MPORT_4_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_0_tile_v_2_MPORT_4_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_0_tile_v_1_MPORT_4_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_0_tile_v_1_MPORT_4_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_0_tile_v_1_MPORT_4_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_0_tile_v_0_MPORT_4_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_0_tile_v_0_MPORT_4_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_0_tile_v_0_MPORT_4_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_1_MPORT_5_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_1_MPORT_5_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_1_MPORT_5_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_0_MPORT_5_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_0_MPORT_5_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_0_MPORT_5_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_0_tile_v_3_MPORT_5_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_0_tile_v_3_MPORT_5_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_0_tile_v_3_MPORT_5_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_0_tile_v_2_MPORT_5_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_0_tile_v_2_MPORT_5_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_0_tile_v_2_MPORT_5_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_0_tile_v_1_MPORT_5_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_0_tile_v_1_MPORT_5_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_0_tile_v_1_MPORT_5_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_0_tile_v_0_MPORT_5_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_0_tile_v_0_MPORT_5_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_0_tile_v_0_MPORT_5_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_0_tile_v_3_MPORT_5_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_0_tile_v_3_MPORT_5_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_0_tile_v_3_MPORT_5_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_0_tile_v_2_MPORT_5_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_0_tile_v_2_MPORT_5_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_0_tile_v_2_MPORT_5_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_0_tile_v_1_MPORT_5_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_0_tile_v_1_MPORT_5_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_0_tile_v_1_MPORT_5_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_0_tile_v_0_MPORT_5_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_0_tile_v_0_MPORT_5_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_0_tile_v_0_MPORT_5_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_1_MPORT_6_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_1_MPORT_6_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_1_MPORT_6_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_0_MPORT_6_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_0_MPORT_6_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_0_MPORT_6_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_0_tile_v_3_MPORT_6_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_0_tile_v_3_MPORT_6_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_0_tile_v_3_MPORT_6_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_0_tile_v_2_MPORT_6_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_0_tile_v_2_MPORT_6_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_0_tile_v_2_MPORT_6_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_0_tile_v_1_MPORT_6_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_0_tile_v_1_MPORT_6_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_0_tile_v_1_MPORT_6_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_0_tile_v_0_MPORT_6_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_0_tile_v_0_MPORT_6_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_0_tile_v_0_MPORT_6_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_0_tile_v_3_MPORT_6_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_0_tile_v_3_MPORT_6_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_0_tile_v_3_MPORT_6_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_0_tile_v_2_MPORT_6_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_0_tile_v_2_MPORT_6_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_0_tile_v_2_MPORT_6_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_0_tile_v_1_MPORT_6_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_0_tile_v_1_MPORT_6_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_0_tile_v_1_MPORT_6_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_0_tile_v_0_MPORT_6_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_0_tile_v_0_MPORT_6_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_0_tile_v_0_MPORT_6_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_3_MPORT_2_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_3_MPORT_2_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_3_MPORT_2_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_2_MPORT_2_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_2_MPORT_2_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_2_MPORT_2_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_1_MPORT_7_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_1_MPORT_7_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_1_MPORT_7_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_0_MPORT_7_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_0_MPORT_7_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_0_MPORT_7_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_0_tile_v_3_MPORT_7_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_0_tile_v_3_MPORT_7_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_0_tile_v_3_MPORT_7_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_0_tile_v_2_MPORT_7_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_0_tile_v_2_MPORT_7_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_0_tile_v_2_MPORT_7_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_0_tile_v_1_MPORT_7_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_0_tile_v_1_MPORT_7_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_0_tile_v_1_MPORT_7_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_0_tile_v_0_MPORT_7_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_0_tile_v_0_MPORT_7_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_0_tile_v_0_MPORT_7_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_0_tile_v_3_MPORT_7_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_0_tile_v_3_MPORT_7_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_0_tile_v_3_MPORT_7_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_0_tile_v_2_MPORT_7_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_0_tile_v_2_MPORT_7_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_0_tile_v_2_MPORT_7_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_0_tile_v_1_MPORT_7_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_0_tile_v_1_MPORT_7_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_0_tile_v_1_MPORT_7_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_0_tile_v_0_MPORT_7_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_0_tile_v_0_MPORT_7_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_0_tile_v_0_MPORT_7_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_1_MPORT_8_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_1_MPORT_8_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_1_MPORT_8_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_0_MPORT_8_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_0_MPORT_8_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_0_MPORT_8_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_0_tile_v_3_MPORT_8_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_0_tile_v_3_MPORT_8_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_0_tile_v_3_MPORT_8_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_0_tile_v_2_MPORT_8_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_0_tile_v_2_MPORT_8_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_0_tile_v_2_MPORT_8_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_0_tile_v_1_MPORT_8_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_0_tile_v_1_MPORT_8_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_0_tile_v_1_MPORT_8_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_0_tile_v_0_MPORT_8_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_0_tile_v_0_MPORT_8_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_0_tile_v_0_MPORT_8_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_0_tile_v_3_MPORT_8_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_0_tile_v_3_MPORT_8_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_0_tile_v_3_MPORT_8_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_0_tile_v_2_MPORT_8_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_0_tile_v_2_MPORT_8_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_0_tile_v_2_MPORT_8_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_0_tile_v_1_MPORT_8_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_0_tile_v_1_MPORT_8_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_0_tile_v_1_MPORT_8_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_0_tile_v_0_MPORT_8_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_0_tile_v_0_MPORT_8_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_0_tile_v_0_MPORT_8_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_3_MPORT_3_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_3_MPORT_3_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_3_MPORT_3_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_2_MPORT_3_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_2_MPORT_3_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_2_MPORT_3_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_1_MPORT_9_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_1_MPORT_9_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_1_MPORT_9_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_0_MPORT_9_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_0_MPORT_9_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_0_MPORT_9_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_0_tile_v_3_MPORT_9_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_0_tile_v_3_MPORT_9_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_0_tile_v_3_MPORT_9_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_0_tile_v_2_MPORT_9_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_0_tile_v_2_MPORT_9_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_0_tile_v_2_MPORT_9_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_0_tile_v_1_MPORT_9_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_0_tile_v_1_MPORT_9_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_0_tile_v_1_MPORT_9_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_0_tile_v_0_MPORT_9_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_0_tile_v_0_MPORT_9_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_0_tile_v_0_MPORT_9_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_0_tile_v_3_MPORT_9_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_0_tile_v_3_MPORT_9_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_0_tile_v_3_MPORT_9_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_0_tile_v_2_MPORT_9_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_0_tile_v_2_MPORT_9_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_0_tile_v_2_MPORT_9_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_0_tile_v_1_MPORT_9_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_0_tile_v_1_MPORT_9_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_0_tile_v_1_MPORT_9_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_0_tile_v_0_MPORT_9_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_0_tile_v_0_MPORT_9_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_0_tile_v_0_MPORT_9_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_1_MPORT_10_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_1_MPORT_10_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_1_MPORT_10_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_0_MPORT_10_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_0_MPORT_10_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_0_MPORT_10_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_0_tile_v_3_MPORT_10_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_0_tile_v_3_MPORT_10_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_0_tile_v_3_MPORT_10_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_0_tile_v_2_MPORT_10_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_0_tile_v_2_MPORT_10_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_0_tile_v_2_MPORT_10_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_0_tile_v_1_MPORT_10_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_0_tile_v_1_MPORT_10_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_0_tile_v_1_MPORT_10_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_0_tile_v_0_MPORT_10_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_0_tile_v_0_MPORT_10_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_0_tile_v_0_MPORT_10_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_0_tile_v_3_MPORT_10_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_0_tile_v_3_MPORT_10_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_0_tile_v_3_MPORT_10_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_0_tile_v_2_MPORT_10_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_0_tile_v_2_MPORT_10_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_0_tile_v_2_MPORT_10_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_0_tile_v_1_MPORT_10_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_0_tile_v_1_MPORT_10_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_0_tile_v_1_MPORT_10_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_0_tile_v_0_MPORT_10_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_0_tile_v_0_MPORT_10_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_0_tile_v_0_MPORT_10_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_1_MPORT_11_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_1_MPORT_11_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_1_MPORT_11_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_0_MPORT_11_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_0_MPORT_11_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_0_MPORT_11_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_0_tile_v_3_MPORT_11_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_0_tile_v_3_MPORT_11_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_0_tile_v_3_MPORT_11_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_0_tile_v_2_MPORT_11_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_0_tile_v_2_MPORT_11_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_0_tile_v_2_MPORT_11_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_0_tile_v_1_MPORT_11_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_0_tile_v_1_MPORT_11_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_0_tile_v_1_MPORT_11_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_0_tile_v_0_MPORT_11_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_0_tile_v_0_MPORT_11_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_0_tile_v_0_MPORT_11_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_0_tile_v_3_MPORT_11_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_0_tile_v_3_MPORT_11_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_0_tile_v_3_MPORT_11_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_0_tile_v_2_MPORT_11_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_0_tile_v_2_MPORT_11_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_0_tile_v_2_MPORT_11_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_0_tile_v_1_MPORT_11_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_0_tile_v_1_MPORT_11_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_0_tile_v_1_MPORT_11_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_0_tile_v_0_MPORT_11_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_0_tile_v_0_MPORT_11_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_0_tile_v_0_MPORT_11_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_1_MPORT_12_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_1_MPORT_12_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_1_MPORT_12_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_0_MPORT_12_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_0_MPORT_12_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_0_MPORT_12_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_0_tile_v_3_MPORT_12_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_0_tile_v_3_MPORT_12_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_0_tile_v_3_MPORT_12_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_0_tile_v_2_MPORT_12_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_0_tile_v_2_MPORT_12_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_0_tile_v_2_MPORT_12_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_0_tile_v_1_MPORT_12_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_0_tile_v_1_MPORT_12_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_0_tile_v_1_MPORT_12_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_0_tile_v_0_MPORT_12_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_0_tile_v_0_MPORT_12_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_0_tile_v_0_MPORT_12_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_0_tile_v_3_MPORT_12_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_0_tile_v_3_MPORT_12_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_0_tile_v_3_MPORT_12_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_0_tile_v_2_MPORT_12_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_0_tile_v_2_MPORT_12_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_0_tile_v_2_MPORT_12_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_0_tile_v_1_MPORT_12_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_0_tile_v_1_MPORT_12_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_0_tile_v_1_MPORT_12_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_0_tile_v_0_MPORT_12_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_0_tile_v_0_MPORT_12_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_0_tile_v_0_MPORT_12_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_3_MPORT_4_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_3_MPORT_4_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_3_MPORT_4_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_2_MPORT_4_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_2_MPORT_4_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_2_MPORT_4_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_1_MPORT_13_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_1_MPORT_13_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_1_MPORT_13_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_0_MPORT_13_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_0_MPORT_13_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_0_MPORT_13_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_0_tile_v_3_MPORT_13_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_0_tile_v_3_MPORT_13_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_0_tile_v_3_MPORT_13_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_0_tile_v_2_MPORT_13_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_0_tile_v_2_MPORT_13_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_0_tile_v_2_MPORT_13_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_0_tile_v_1_MPORT_13_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_0_tile_v_1_MPORT_13_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_0_tile_v_1_MPORT_13_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_0_tile_v_0_MPORT_13_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_0_tile_v_0_MPORT_13_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_0_tile_v_0_MPORT_13_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_0_tile_v_3_MPORT_13_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_0_tile_v_3_MPORT_13_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_0_tile_v_3_MPORT_13_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_0_tile_v_2_MPORT_13_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_0_tile_v_2_MPORT_13_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_0_tile_v_2_MPORT_13_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_0_tile_v_1_MPORT_13_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_0_tile_v_1_MPORT_13_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_0_tile_v_1_MPORT_13_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_0_tile_v_0_MPORT_13_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_0_tile_v_0_MPORT_13_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_0_tile_v_0_MPORT_13_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_1_MPORT_14_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_1_MPORT_14_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_1_MPORT_14_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_0_MPORT_14_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_0_MPORT_14_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_0_MPORT_14_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_0_tile_v_3_MPORT_14_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_0_tile_v_3_MPORT_14_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_0_tile_v_3_MPORT_14_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_0_tile_v_2_MPORT_14_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_0_tile_v_2_MPORT_14_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_0_tile_v_2_MPORT_14_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_0_tile_v_1_MPORT_14_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_0_tile_v_1_MPORT_14_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_0_tile_v_1_MPORT_14_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_0_tile_v_0_MPORT_14_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_0_tile_v_0_MPORT_14_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_0_tile_v_0_MPORT_14_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_0_tile_v_3_MPORT_14_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_0_tile_v_3_MPORT_14_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_0_tile_v_3_MPORT_14_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_0_tile_v_2_MPORT_14_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_0_tile_v_2_MPORT_14_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_0_tile_v_2_MPORT_14_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_0_tile_v_1_MPORT_14_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_0_tile_v_1_MPORT_14_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_0_tile_v_1_MPORT_14_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_0_tile_v_0_MPORT_14_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_0_tile_v_0_MPORT_14_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_0_tile_v_0_MPORT_14_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_3_MPORT_5_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_3_MPORT_5_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_3_MPORT_5_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_2_MPORT_5_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_2_MPORT_5_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_2_MPORT_5_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_1_MPORT_15_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_1_MPORT_15_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_1_MPORT_15_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_0_MPORT_15_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_0_MPORT_15_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_0_MPORT_15_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_0_tile_v_3_MPORT_15_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_0_tile_v_3_MPORT_15_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_0_tile_v_3_MPORT_15_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_0_tile_v_2_MPORT_15_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_0_tile_v_2_MPORT_15_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_0_tile_v_2_MPORT_15_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_0_tile_v_1_MPORT_15_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_0_tile_v_1_MPORT_15_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_0_tile_v_1_MPORT_15_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_0_tile_v_0_MPORT_15_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_0_tile_v_0_MPORT_15_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_0_tile_v_0_MPORT_15_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_0_tile_v_3_MPORT_15_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_0_tile_v_3_MPORT_15_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_0_tile_v_3_MPORT_15_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_0_tile_v_2_MPORT_15_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_0_tile_v_2_MPORT_15_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_0_tile_v_2_MPORT_15_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_0_tile_v_1_MPORT_15_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_0_tile_v_1_MPORT_15_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_0_tile_v_1_MPORT_15_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_0_tile_v_0_MPORT_15_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_0_tile_v_0_MPORT_15_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_0_tile_v_0_MPORT_15_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_1_MPORT_16_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_1_MPORT_16_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_1_MPORT_16_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_0_MPORT_16_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_0_MPORT_16_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_0_MPORT_16_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_0_tile_v_3_MPORT_16_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_0_tile_v_3_MPORT_16_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_0_tile_v_3_MPORT_16_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_0_tile_v_2_MPORT_16_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_0_tile_v_2_MPORT_16_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_0_tile_v_2_MPORT_16_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_0_tile_v_1_MPORT_16_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_0_tile_v_1_MPORT_16_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_0_tile_v_1_MPORT_16_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_0_tile_v_0_MPORT_16_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_0_tile_v_0_MPORT_16_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_0_tile_v_0_MPORT_16_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_0_tile_v_3_MPORT_16_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_0_tile_v_3_MPORT_16_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_0_tile_v_3_MPORT_16_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_0_tile_v_2_MPORT_16_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_0_tile_v_2_MPORT_16_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_0_tile_v_2_MPORT_16_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_0_tile_v_1_MPORT_16_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_0_tile_v_1_MPORT_16_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_0_tile_v_1_MPORT_16_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_0_tile_v_0_MPORT_16_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_0_tile_v_0_MPORT_16_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_0_tile_v_0_MPORT_16_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_1_MPORT_17_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_1_MPORT_17_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_1_MPORT_17_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_0_MPORT_17_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_0_MPORT_17_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_0_MPORT_17_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_0_tile_v_3_MPORT_17_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_0_tile_v_3_MPORT_17_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_0_tile_v_3_MPORT_17_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_0_tile_v_2_MPORT_17_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_0_tile_v_2_MPORT_17_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_0_tile_v_2_MPORT_17_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_0_tile_v_1_MPORT_17_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_0_tile_v_1_MPORT_17_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_0_tile_v_1_MPORT_17_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_0_tile_v_0_MPORT_17_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_0_tile_v_0_MPORT_17_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_0_tile_v_0_MPORT_17_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_0_tile_v_3_MPORT_17_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_0_tile_v_3_MPORT_17_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_0_tile_v_3_MPORT_17_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_0_tile_v_2_MPORT_17_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_0_tile_v_2_MPORT_17_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_0_tile_v_2_MPORT_17_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_0_tile_v_1_MPORT_17_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_0_tile_v_1_MPORT_17_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_0_tile_v_1_MPORT_17_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_0_tile_v_0_MPORT_17_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_0_tile_v_0_MPORT_17_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_0_tile_v_0_MPORT_17_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_1_MPORT_18_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_1_MPORT_18_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_1_MPORT_18_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_0_MPORT_18_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_0_MPORT_18_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_0_MPORT_18_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_0_tile_v_3_MPORT_18_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_0_tile_v_3_MPORT_18_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_0_tile_v_3_MPORT_18_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_0_tile_v_2_MPORT_18_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_0_tile_v_2_MPORT_18_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_0_tile_v_2_MPORT_18_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_0_tile_v_1_MPORT_18_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_0_tile_v_1_MPORT_18_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_0_tile_v_1_MPORT_18_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_0_tile_v_0_MPORT_18_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_0_tile_v_0_MPORT_18_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_0_tile_v_0_MPORT_18_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_0_tile_v_3_MPORT_18_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_0_tile_v_3_MPORT_18_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_0_tile_v_3_MPORT_18_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_0_tile_v_2_MPORT_18_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_0_tile_v_2_MPORT_18_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_0_tile_v_2_MPORT_18_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_0_tile_v_1_MPORT_18_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_0_tile_v_1_MPORT_18_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_0_tile_v_1_MPORT_18_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_0_tile_v_0_MPORT_18_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_0_tile_v_0_MPORT_18_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_0_tile_v_0_MPORT_18_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_3_MPORT_6_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_3_MPORT_6_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_3_MPORT_6_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_2_MPORT_6_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_2_MPORT_6_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_2_MPORT_6_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_1_MPORT_19_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_1_MPORT_19_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_1_MPORT_19_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_0_MPORT_19_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_0_MPORT_19_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_0_MPORT_19_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_0_tile_v_3_MPORT_19_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_0_tile_v_3_MPORT_19_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_0_tile_v_3_MPORT_19_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_0_tile_v_2_MPORT_19_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_0_tile_v_2_MPORT_19_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_0_tile_v_2_MPORT_19_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_0_tile_v_1_MPORT_19_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_0_tile_v_1_MPORT_19_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_0_tile_v_1_MPORT_19_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_0_tile_v_0_MPORT_19_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_0_tile_v_0_MPORT_19_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_0_tile_v_0_MPORT_19_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_0_tile_v_3_MPORT_19_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_0_tile_v_3_MPORT_19_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_0_tile_v_3_MPORT_19_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_0_tile_v_2_MPORT_19_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_0_tile_v_2_MPORT_19_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_0_tile_v_2_MPORT_19_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_0_tile_v_1_MPORT_19_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_0_tile_v_1_MPORT_19_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_0_tile_v_1_MPORT_19_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_0_tile_v_0_MPORT_19_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_0_tile_v_0_MPORT_19_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_0_tile_v_0_MPORT_19_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_1_MPORT_20_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_1_MPORT_20_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_1_MPORT_20_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_0_MPORT_20_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_0_MPORT_20_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_0_MPORT_20_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_0_tile_v_3_MPORT_20_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_0_tile_v_3_MPORT_20_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_0_tile_v_3_MPORT_20_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_0_tile_v_2_MPORT_20_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_0_tile_v_2_MPORT_20_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_0_tile_v_2_MPORT_20_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_0_tile_v_1_MPORT_20_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_0_tile_v_1_MPORT_20_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_0_tile_v_1_MPORT_20_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_0_tile_v_0_MPORT_20_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_0_tile_v_0_MPORT_20_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_0_tile_v_0_MPORT_20_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_0_tile_v_3_MPORT_20_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_0_tile_v_3_MPORT_20_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_0_tile_v_3_MPORT_20_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_0_tile_v_2_MPORT_20_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_0_tile_v_2_MPORT_20_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_0_tile_v_2_MPORT_20_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_0_tile_v_1_MPORT_20_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_0_tile_v_1_MPORT_20_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_0_tile_v_1_MPORT_20_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_0_tile_v_0_MPORT_20_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_0_tile_v_0_MPORT_20_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_0_tile_v_0_MPORT_20_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_3_MPORT_7_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_3_MPORT_7_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_3_MPORT_7_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_2_MPORT_7_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_2_MPORT_7_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_2_MPORT_7_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_1_MPORT_21_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_1_MPORT_21_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_1_MPORT_21_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_0_MPORT_21_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_0_MPORT_21_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_0_MPORT_21_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_0_tile_v_3_MPORT_21_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_0_tile_v_3_MPORT_21_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_0_tile_v_3_MPORT_21_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_0_tile_v_2_MPORT_21_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_0_tile_v_2_MPORT_21_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_0_tile_v_2_MPORT_21_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_0_tile_v_1_MPORT_21_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_0_tile_v_1_MPORT_21_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_0_tile_v_1_MPORT_21_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_0_tile_v_0_MPORT_21_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_0_tile_v_0_MPORT_21_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_0_tile_v_0_MPORT_21_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_0_tile_v_3_MPORT_21_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_0_tile_v_3_MPORT_21_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_0_tile_v_3_MPORT_21_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_0_tile_v_2_MPORT_21_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_0_tile_v_2_MPORT_21_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_0_tile_v_2_MPORT_21_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_0_tile_v_1_MPORT_21_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_0_tile_v_1_MPORT_21_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_0_tile_v_1_MPORT_21_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_0_tile_v_0_MPORT_21_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_0_tile_v_0_MPORT_21_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_0_tile_v_0_MPORT_21_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_1_MPORT_22_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_1_MPORT_22_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_1_MPORT_22_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_0_MPORT_22_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_0_MPORT_22_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_0_MPORT_22_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_0_tile_v_3_MPORT_22_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_0_tile_v_3_MPORT_22_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_0_tile_v_3_MPORT_22_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_0_tile_v_2_MPORT_22_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_0_tile_v_2_MPORT_22_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_0_tile_v_2_MPORT_22_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_0_tile_v_1_MPORT_22_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_0_tile_v_1_MPORT_22_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_0_tile_v_1_MPORT_22_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_0_tile_v_0_MPORT_22_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_0_tile_v_0_MPORT_22_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_0_tile_v_0_MPORT_22_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_0_tile_v_3_MPORT_22_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_0_tile_v_3_MPORT_22_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_0_tile_v_3_MPORT_22_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_0_tile_v_2_MPORT_22_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_0_tile_v_2_MPORT_22_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_0_tile_v_2_MPORT_22_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_0_tile_v_1_MPORT_22_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_0_tile_v_1_MPORT_22_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_0_tile_v_1_MPORT_22_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_0_tile_v_0_MPORT_22_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_0_tile_v_0_MPORT_22_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_0_tile_v_0_MPORT_22_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_1_MPORT_23_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_1_MPORT_23_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_1_MPORT_23_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_0_MPORT_23_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_0_MPORT_23_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_0_MPORT_23_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_0_tile_v_3_MPORT_23_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_0_tile_v_3_MPORT_23_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_0_tile_v_3_MPORT_23_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_0_tile_v_2_MPORT_23_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_0_tile_v_2_MPORT_23_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_0_tile_v_2_MPORT_23_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_0_tile_v_1_MPORT_23_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_0_tile_v_1_MPORT_23_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_0_tile_v_1_MPORT_23_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_0_tile_v_0_MPORT_23_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_0_tile_v_0_MPORT_23_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_0_tile_v_0_MPORT_23_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_0_tile_v_3_MPORT_23_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_0_tile_v_3_MPORT_23_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_0_tile_v_3_MPORT_23_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_0_tile_v_2_MPORT_23_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_0_tile_v_2_MPORT_23_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_0_tile_v_2_MPORT_23_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_0_tile_v_1_MPORT_23_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_0_tile_v_1_MPORT_23_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_0_tile_v_1_MPORT_23_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_0_tile_v_0_MPORT_23_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_0_tile_v_0_MPORT_23_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_0_tile_v_0_MPORT_23_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_1_MPORT_24_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_1_MPORT_24_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_1_MPORT_24_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_0_MPORT_24_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_0_MPORT_24_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_0_MPORT_24_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_1_tile_v_3_MPORT_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_1_tile_v_3_MPORT_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_1_tile_v_3_MPORT_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_1_tile_v_2_MPORT_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_1_tile_v_2_MPORT_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_1_tile_v_2_MPORT_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_1_tile_v_1_MPORT_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_1_tile_v_1_MPORT_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_1_tile_v_1_MPORT_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_1_tile_v_0_MPORT_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_1_tile_v_0_MPORT_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_1_tile_v_0_MPORT_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_1_tile_v_3_MPORT_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_1_tile_v_3_MPORT_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_1_tile_v_3_MPORT_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_1_tile_v_2_MPORT_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_1_tile_v_2_MPORT_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_1_tile_v_2_MPORT_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_1_tile_v_1_MPORT_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_1_tile_v_1_MPORT_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_1_tile_v_1_MPORT_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_1_tile_v_0_MPORT_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_1_tile_v_0_MPORT_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_1_tile_v_0_MPORT_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_3_MPORT_8_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_3_MPORT_8_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_3_MPORT_8_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_2_MPORT_8_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_2_MPORT_8_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_2_MPORT_8_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_1_MPORT_25_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_1_MPORT_25_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_1_MPORT_25_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_0_MPORT_25_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_0_MPORT_25_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_0_MPORT_25_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_1_tile_v_3_MPORT_1_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_1_tile_v_3_MPORT_1_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_1_tile_v_3_MPORT_1_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_1_tile_v_2_MPORT_1_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_1_tile_v_2_MPORT_1_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_1_tile_v_2_MPORT_1_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_1_tile_v_1_MPORT_1_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_1_tile_v_1_MPORT_1_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_1_tile_v_1_MPORT_1_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_1_tile_v_0_MPORT_1_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_1_tile_v_0_MPORT_1_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_1_tile_v_0_MPORT_1_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_1_tile_v_3_MPORT_1_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_1_tile_v_3_MPORT_1_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_1_tile_v_3_MPORT_1_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_1_tile_v_2_MPORT_1_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_1_tile_v_2_MPORT_1_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_1_tile_v_2_MPORT_1_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_1_tile_v_1_MPORT_1_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_1_tile_v_1_MPORT_1_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_1_tile_v_1_MPORT_1_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_1_tile_v_0_MPORT_1_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_1_tile_v_0_MPORT_1_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_1_tile_v_0_MPORT_1_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_1_MPORT_26_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_1_MPORT_26_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_1_MPORT_26_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_0_MPORT_26_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_0_MPORT_26_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_0_MPORT_26_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_1_tile_v_3_MPORT_2_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_1_tile_v_3_MPORT_2_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_1_tile_v_3_MPORT_2_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_1_tile_v_2_MPORT_2_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_1_tile_v_2_MPORT_2_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_1_tile_v_2_MPORT_2_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_1_tile_v_1_MPORT_2_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_1_tile_v_1_MPORT_2_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_1_tile_v_1_MPORT_2_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_1_tile_v_0_MPORT_2_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_1_tile_v_0_MPORT_2_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_1_tile_v_0_MPORT_2_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_1_tile_v_3_MPORT_2_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_1_tile_v_3_MPORT_2_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_1_tile_v_3_MPORT_2_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_1_tile_v_2_MPORT_2_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_1_tile_v_2_MPORT_2_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_1_tile_v_2_MPORT_2_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_1_tile_v_1_MPORT_2_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_1_tile_v_1_MPORT_2_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_1_tile_v_1_MPORT_2_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_1_tile_v_0_MPORT_2_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_1_tile_v_0_MPORT_2_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_1_tile_v_0_MPORT_2_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_3_MPORT_9_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_3_MPORT_9_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_3_MPORT_9_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_2_MPORT_9_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_2_MPORT_9_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_2_MPORT_9_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_1_MPORT_27_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_1_MPORT_27_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_1_MPORT_27_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_0_MPORT_27_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_0_MPORT_27_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_0_MPORT_27_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_1_tile_v_3_MPORT_3_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_1_tile_v_3_MPORT_3_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_1_tile_v_3_MPORT_3_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_1_tile_v_2_MPORT_3_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_1_tile_v_2_MPORT_3_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_1_tile_v_2_MPORT_3_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_1_tile_v_1_MPORT_3_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_1_tile_v_1_MPORT_3_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_1_tile_v_1_MPORT_3_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_1_tile_v_0_MPORT_3_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_1_tile_v_0_MPORT_3_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_1_tile_v_0_MPORT_3_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_1_tile_v_3_MPORT_3_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_1_tile_v_3_MPORT_3_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_1_tile_v_3_MPORT_3_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_1_tile_v_2_MPORT_3_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_1_tile_v_2_MPORT_3_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_1_tile_v_2_MPORT_3_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_1_tile_v_1_MPORT_3_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_1_tile_v_1_MPORT_3_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_1_tile_v_1_MPORT_3_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_1_tile_v_0_MPORT_3_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_1_tile_v_0_MPORT_3_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_1_tile_v_0_MPORT_3_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_1_MPORT_28_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_1_MPORT_28_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_1_MPORT_28_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_0_MPORT_28_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_0_MPORT_28_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_0_MPORT_28_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_1_tile_v_3_MPORT_4_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_1_tile_v_3_MPORT_4_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_1_tile_v_3_MPORT_4_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_1_tile_v_2_MPORT_4_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_1_tile_v_2_MPORT_4_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_1_tile_v_2_MPORT_4_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_1_tile_v_1_MPORT_4_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_1_tile_v_1_MPORT_4_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_1_tile_v_1_MPORT_4_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_1_tile_v_0_MPORT_4_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_1_tile_v_0_MPORT_4_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_1_tile_v_0_MPORT_4_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_1_tile_v_3_MPORT_4_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_1_tile_v_3_MPORT_4_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_1_tile_v_3_MPORT_4_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_1_tile_v_2_MPORT_4_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_1_tile_v_2_MPORT_4_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_1_tile_v_2_MPORT_4_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_1_tile_v_1_MPORT_4_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_1_tile_v_1_MPORT_4_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_1_tile_v_1_MPORT_4_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_1_tile_v_0_MPORT_4_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_1_tile_v_0_MPORT_4_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_1_tile_v_0_MPORT_4_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_1_MPORT_29_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_1_MPORT_29_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_1_MPORT_29_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_0_MPORT_29_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_0_MPORT_29_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_0_MPORT_29_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_1_tile_v_3_MPORT_5_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_1_tile_v_3_MPORT_5_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_1_tile_v_3_MPORT_5_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_1_tile_v_2_MPORT_5_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_1_tile_v_2_MPORT_5_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_1_tile_v_2_MPORT_5_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_1_tile_v_1_MPORT_5_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_1_tile_v_1_MPORT_5_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_1_tile_v_1_MPORT_5_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_1_tile_v_0_MPORT_5_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_1_tile_v_0_MPORT_5_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_1_tile_v_0_MPORT_5_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_1_tile_v_3_MPORT_5_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_1_tile_v_3_MPORT_5_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_1_tile_v_3_MPORT_5_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_1_tile_v_2_MPORT_5_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_1_tile_v_2_MPORT_5_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_1_tile_v_2_MPORT_5_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_1_tile_v_1_MPORT_5_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_1_tile_v_1_MPORT_5_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_1_tile_v_1_MPORT_5_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_1_tile_v_0_MPORT_5_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_1_tile_v_0_MPORT_5_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_1_tile_v_0_MPORT_5_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_1_MPORT_30_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_1_MPORT_30_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_1_MPORT_30_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_0_MPORT_30_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_0_MPORT_30_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_0_MPORT_30_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_1_tile_v_3_MPORT_6_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_1_tile_v_3_MPORT_6_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_1_tile_v_3_MPORT_6_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_1_tile_v_2_MPORT_6_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_1_tile_v_2_MPORT_6_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_1_tile_v_2_MPORT_6_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_1_tile_v_1_MPORT_6_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_1_tile_v_1_MPORT_6_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_1_tile_v_1_MPORT_6_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_1_tile_v_0_MPORT_6_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_1_tile_v_0_MPORT_6_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_1_tile_v_0_MPORT_6_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_1_tile_v_3_MPORT_6_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_1_tile_v_3_MPORT_6_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_1_tile_v_3_MPORT_6_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_1_tile_v_2_MPORT_6_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_1_tile_v_2_MPORT_6_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_1_tile_v_2_MPORT_6_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_1_tile_v_1_MPORT_6_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_1_tile_v_1_MPORT_6_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_1_tile_v_1_MPORT_6_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_1_tile_v_0_MPORT_6_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_1_tile_v_0_MPORT_6_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_1_tile_v_0_MPORT_6_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_3_MPORT_10_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_3_MPORT_10_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_3_MPORT_10_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_2_MPORT_10_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_2_MPORT_10_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_2_MPORT_10_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_1_MPORT_31_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_1_MPORT_31_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_1_MPORT_31_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_0_MPORT_31_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_0_MPORT_31_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_0_MPORT_31_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_1_tile_v_3_MPORT_7_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_1_tile_v_3_MPORT_7_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_1_tile_v_3_MPORT_7_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_1_tile_v_2_MPORT_7_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_1_tile_v_2_MPORT_7_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_1_tile_v_2_MPORT_7_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_1_tile_v_1_MPORT_7_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_1_tile_v_1_MPORT_7_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_1_tile_v_1_MPORT_7_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_1_tile_v_0_MPORT_7_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_1_tile_v_0_MPORT_7_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_1_tile_v_0_MPORT_7_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_1_tile_v_3_MPORT_7_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_1_tile_v_3_MPORT_7_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_1_tile_v_3_MPORT_7_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_1_tile_v_2_MPORT_7_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_1_tile_v_2_MPORT_7_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_1_tile_v_2_MPORT_7_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_1_tile_v_1_MPORT_7_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_1_tile_v_1_MPORT_7_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_1_tile_v_1_MPORT_7_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_1_tile_v_0_MPORT_7_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_1_tile_v_0_MPORT_7_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_1_tile_v_0_MPORT_7_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_1_MPORT_32_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_1_MPORT_32_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_1_MPORT_32_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_0_MPORT_32_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_0_MPORT_32_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_0_MPORT_32_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_1_tile_v_3_MPORT_8_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_1_tile_v_3_MPORT_8_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_1_tile_v_3_MPORT_8_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_1_tile_v_2_MPORT_8_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_1_tile_v_2_MPORT_8_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_1_tile_v_2_MPORT_8_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_1_tile_v_1_MPORT_8_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_1_tile_v_1_MPORT_8_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_1_tile_v_1_MPORT_8_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_1_tile_v_0_MPORT_8_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_1_tile_v_0_MPORT_8_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_1_tile_v_0_MPORT_8_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_1_tile_v_3_MPORT_8_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_1_tile_v_3_MPORT_8_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_1_tile_v_3_MPORT_8_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_1_tile_v_2_MPORT_8_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_1_tile_v_2_MPORT_8_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_1_tile_v_2_MPORT_8_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_1_tile_v_1_MPORT_8_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_1_tile_v_1_MPORT_8_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_1_tile_v_1_MPORT_8_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_1_tile_v_0_MPORT_8_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_1_tile_v_0_MPORT_8_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_1_tile_v_0_MPORT_8_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_3_MPORT_11_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_3_MPORT_11_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_3_MPORT_11_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_2_MPORT_11_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_2_MPORT_11_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_2_MPORT_11_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_1_MPORT_33_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_1_MPORT_33_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_1_MPORT_33_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_0_MPORT_33_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_0_MPORT_33_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_0_MPORT_33_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_1_tile_v_3_MPORT_9_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_1_tile_v_3_MPORT_9_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_1_tile_v_3_MPORT_9_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_1_tile_v_2_MPORT_9_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_1_tile_v_2_MPORT_9_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_1_tile_v_2_MPORT_9_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_1_tile_v_1_MPORT_9_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_1_tile_v_1_MPORT_9_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_1_tile_v_1_MPORT_9_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_1_tile_v_0_MPORT_9_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_1_tile_v_0_MPORT_9_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_1_tile_v_0_MPORT_9_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_1_tile_v_3_MPORT_9_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_1_tile_v_3_MPORT_9_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_1_tile_v_3_MPORT_9_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_1_tile_v_2_MPORT_9_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_1_tile_v_2_MPORT_9_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_1_tile_v_2_MPORT_9_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_1_tile_v_1_MPORT_9_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_1_tile_v_1_MPORT_9_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_1_tile_v_1_MPORT_9_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_1_tile_v_0_MPORT_9_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_1_tile_v_0_MPORT_9_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_1_tile_v_0_MPORT_9_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_1_MPORT_34_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_1_MPORT_34_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_1_MPORT_34_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_0_MPORT_34_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_0_MPORT_34_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_0_MPORT_34_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_1_tile_v_3_MPORT_10_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_1_tile_v_3_MPORT_10_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_1_tile_v_3_MPORT_10_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_1_tile_v_2_MPORT_10_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_1_tile_v_2_MPORT_10_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_1_tile_v_2_MPORT_10_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_1_tile_v_1_MPORT_10_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_1_tile_v_1_MPORT_10_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_1_tile_v_1_MPORT_10_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_1_tile_v_0_MPORT_10_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_1_tile_v_0_MPORT_10_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_1_tile_v_0_MPORT_10_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_1_tile_v_3_MPORT_10_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_1_tile_v_3_MPORT_10_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_1_tile_v_3_MPORT_10_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_1_tile_v_2_MPORT_10_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_1_tile_v_2_MPORT_10_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_1_tile_v_2_MPORT_10_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_1_tile_v_1_MPORT_10_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_1_tile_v_1_MPORT_10_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_1_tile_v_1_MPORT_10_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_1_tile_v_0_MPORT_10_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_1_tile_v_0_MPORT_10_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_1_tile_v_0_MPORT_10_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_1_MPORT_35_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_1_MPORT_35_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_1_MPORT_35_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_0_MPORT_35_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_0_MPORT_35_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_0_MPORT_35_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_1_tile_v_3_MPORT_11_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_1_tile_v_3_MPORT_11_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_1_tile_v_3_MPORT_11_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_1_tile_v_2_MPORT_11_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_1_tile_v_2_MPORT_11_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_1_tile_v_2_MPORT_11_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_1_tile_v_1_MPORT_11_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_1_tile_v_1_MPORT_11_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_1_tile_v_1_MPORT_11_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_1_tile_v_0_MPORT_11_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_1_tile_v_0_MPORT_11_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_1_tile_v_0_MPORT_11_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_1_tile_v_3_MPORT_11_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_1_tile_v_3_MPORT_11_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_1_tile_v_3_MPORT_11_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_1_tile_v_2_MPORT_11_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_1_tile_v_2_MPORT_11_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_1_tile_v_2_MPORT_11_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_1_tile_v_1_MPORT_11_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_1_tile_v_1_MPORT_11_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_1_tile_v_1_MPORT_11_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_1_tile_v_0_MPORT_11_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_1_tile_v_0_MPORT_11_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_1_tile_v_0_MPORT_11_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_1_MPORT_36_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_1_MPORT_36_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_1_MPORT_36_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_0_MPORT_36_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_0_MPORT_36_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_0_MPORT_36_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_1_tile_v_3_MPORT_12_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_1_tile_v_3_MPORT_12_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_1_tile_v_3_MPORT_12_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_1_tile_v_2_MPORT_12_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_1_tile_v_2_MPORT_12_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_1_tile_v_2_MPORT_12_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_1_tile_v_1_MPORT_12_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_1_tile_v_1_MPORT_12_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_1_tile_v_1_MPORT_12_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_1_tile_v_0_MPORT_12_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_1_tile_v_0_MPORT_12_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_1_tile_v_0_MPORT_12_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_1_tile_v_3_MPORT_12_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_1_tile_v_3_MPORT_12_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_1_tile_v_3_MPORT_12_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_1_tile_v_2_MPORT_12_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_1_tile_v_2_MPORT_12_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_1_tile_v_2_MPORT_12_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_1_tile_v_1_MPORT_12_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_1_tile_v_1_MPORT_12_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_1_tile_v_1_MPORT_12_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_1_tile_v_0_MPORT_12_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_1_tile_v_0_MPORT_12_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_1_tile_v_0_MPORT_12_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_3_MPORT_12_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_3_MPORT_12_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_3_MPORT_12_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_2_MPORT_12_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_2_MPORT_12_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_2_MPORT_12_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_1_MPORT_37_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_1_MPORT_37_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_1_MPORT_37_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_0_MPORT_37_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_0_MPORT_37_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_0_MPORT_37_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_1_tile_v_3_MPORT_13_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_1_tile_v_3_MPORT_13_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_1_tile_v_3_MPORT_13_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_1_tile_v_2_MPORT_13_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_1_tile_v_2_MPORT_13_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_1_tile_v_2_MPORT_13_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_1_tile_v_1_MPORT_13_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_1_tile_v_1_MPORT_13_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_1_tile_v_1_MPORT_13_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_1_tile_v_0_MPORT_13_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_1_tile_v_0_MPORT_13_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_1_tile_v_0_MPORT_13_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_1_tile_v_3_MPORT_13_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_1_tile_v_3_MPORT_13_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_1_tile_v_3_MPORT_13_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_1_tile_v_2_MPORT_13_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_1_tile_v_2_MPORT_13_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_1_tile_v_2_MPORT_13_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_1_tile_v_1_MPORT_13_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_1_tile_v_1_MPORT_13_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_1_tile_v_1_MPORT_13_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_1_tile_v_0_MPORT_13_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_1_tile_v_0_MPORT_13_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_1_tile_v_0_MPORT_13_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_1_MPORT_38_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_1_MPORT_38_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_1_MPORT_38_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_0_MPORT_38_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_0_MPORT_38_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_0_MPORT_38_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_1_tile_v_3_MPORT_14_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_1_tile_v_3_MPORT_14_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_1_tile_v_3_MPORT_14_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_1_tile_v_2_MPORT_14_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_1_tile_v_2_MPORT_14_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_1_tile_v_2_MPORT_14_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_1_tile_v_1_MPORT_14_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_1_tile_v_1_MPORT_14_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_1_tile_v_1_MPORT_14_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_1_tile_v_0_MPORT_14_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_1_tile_v_0_MPORT_14_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_1_tile_v_0_MPORT_14_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_1_tile_v_3_MPORT_14_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_1_tile_v_3_MPORT_14_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_1_tile_v_3_MPORT_14_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_1_tile_v_2_MPORT_14_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_1_tile_v_2_MPORT_14_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_1_tile_v_2_MPORT_14_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_1_tile_v_1_MPORT_14_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_1_tile_v_1_MPORT_14_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_1_tile_v_1_MPORT_14_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_1_tile_v_0_MPORT_14_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_1_tile_v_0_MPORT_14_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_1_tile_v_0_MPORT_14_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_3_MPORT_13_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_3_MPORT_13_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_3_MPORT_13_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_2_MPORT_13_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_2_MPORT_13_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_2_MPORT_13_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_1_MPORT_39_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_1_MPORT_39_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_1_MPORT_39_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_0_MPORT_39_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_0_MPORT_39_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_0_MPORT_39_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_1_tile_v_3_MPORT_15_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_1_tile_v_3_MPORT_15_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_1_tile_v_3_MPORT_15_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_1_tile_v_2_MPORT_15_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_1_tile_v_2_MPORT_15_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_1_tile_v_2_MPORT_15_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_1_tile_v_1_MPORT_15_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_1_tile_v_1_MPORT_15_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_1_tile_v_1_MPORT_15_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_1_tile_v_0_MPORT_15_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_1_tile_v_0_MPORT_15_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_1_tile_v_0_MPORT_15_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_1_tile_v_3_MPORT_15_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_1_tile_v_3_MPORT_15_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_1_tile_v_3_MPORT_15_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_1_tile_v_2_MPORT_15_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_1_tile_v_2_MPORT_15_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_1_tile_v_2_MPORT_15_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_1_tile_v_1_MPORT_15_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_1_tile_v_1_MPORT_15_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_1_tile_v_1_MPORT_15_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_1_tile_v_0_MPORT_15_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_1_tile_v_0_MPORT_15_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_1_tile_v_0_MPORT_15_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_1_MPORT_40_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_1_MPORT_40_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_1_MPORT_40_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_0_MPORT_40_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_0_MPORT_40_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_0_MPORT_40_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_1_tile_v_3_MPORT_16_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_1_tile_v_3_MPORT_16_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_1_tile_v_3_MPORT_16_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_1_tile_v_2_MPORT_16_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_1_tile_v_2_MPORT_16_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_1_tile_v_2_MPORT_16_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_1_tile_v_1_MPORT_16_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_1_tile_v_1_MPORT_16_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_1_tile_v_1_MPORT_16_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_1_tile_v_0_MPORT_16_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_1_tile_v_0_MPORT_16_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_1_tile_v_0_MPORT_16_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_1_tile_v_3_MPORT_16_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_1_tile_v_3_MPORT_16_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_1_tile_v_3_MPORT_16_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_1_tile_v_2_MPORT_16_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_1_tile_v_2_MPORT_16_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_1_tile_v_2_MPORT_16_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_1_tile_v_1_MPORT_16_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_1_tile_v_1_MPORT_16_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_1_tile_v_1_MPORT_16_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_1_tile_v_0_MPORT_16_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_1_tile_v_0_MPORT_16_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_1_tile_v_0_MPORT_16_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_1_MPORT_41_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_1_MPORT_41_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_1_MPORT_41_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_0_MPORT_41_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_0_MPORT_41_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_0_MPORT_41_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_1_tile_v_3_MPORT_17_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_1_tile_v_3_MPORT_17_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_1_tile_v_3_MPORT_17_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_1_tile_v_2_MPORT_17_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_1_tile_v_2_MPORT_17_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_1_tile_v_2_MPORT_17_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_1_tile_v_1_MPORT_17_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_1_tile_v_1_MPORT_17_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_1_tile_v_1_MPORT_17_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_1_tile_v_0_MPORT_17_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_1_tile_v_0_MPORT_17_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_1_tile_v_0_MPORT_17_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_1_tile_v_3_MPORT_17_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_1_tile_v_3_MPORT_17_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_1_tile_v_3_MPORT_17_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_1_tile_v_2_MPORT_17_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_1_tile_v_2_MPORT_17_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_1_tile_v_2_MPORT_17_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_1_tile_v_1_MPORT_17_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_1_tile_v_1_MPORT_17_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_1_tile_v_1_MPORT_17_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_1_tile_v_0_MPORT_17_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_1_tile_v_0_MPORT_17_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_1_tile_v_0_MPORT_17_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_1_MPORT_42_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_1_MPORT_42_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_1_MPORT_42_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_0_MPORT_42_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_0_MPORT_42_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_0_MPORT_42_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_1_tile_v_3_MPORT_18_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_1_tile_v_3_MPORT_18_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_1_tile_v_3_MPORT_18_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_1_tile_v_2_MPORT_18_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_1_tile_v_2_MPORT_18_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_1_tile_v_2_MPORT_18_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_1_tile_v_1_MPORT_18_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_1_tile_v_1_MPORT_18_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_1_tile_v_1_MPORT_18_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_1_tile_v_0_MPORT_18_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_1_tile_v_0_MPORT_18_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_1_tile_v_0_MPORT_18_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_1_tile_v_3_MPORT_18_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_1_tile_v_3_MPORT_18_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_1_tile_v_3_MPORT_18_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_1_tile_v_2_MPORT_18_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_1_tile_v_2_MPORT_18_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_1_tile_v_2_MPORT_18_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_1_tile_v_1_MPORT_18_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_1_tile_v_1_MPORT_18_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_1_tile_v_1_MPORT_18_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_1_tile_v_0_MPORT_18_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_1_tile_v_0_MPORT_18_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_1_tile_v_0_MPORT_18_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_3_MPORT_14_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_3_MPORT_14_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_3_MPORT_14_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_2_MPORT_14_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_2_MPORT_14_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_2_MPORT_14_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_1_MPORT_43_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_1_MPORT_43_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_1_MPORT_43_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_0_MPORT_43_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_0_MPORT_43_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_0_MPORT_43_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_1_tile_v_3_MPORT_19_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_1_tile_v_3_MPORT_19_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_1_tile_v_3_MPORT_19_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_1_tile_v_2_MPORT_19_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_1_tile_v_2_MPORT_19_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_1_tile_v_2_MPORT_19_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_1_tile_v_1_MPORT_19_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_1_tile_v_1_MPORT_19_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_1_tile_v_1_MPORT_19_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_1_tile_v_0_MPORT_19_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_1_tile_v_0_MPORT_19_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_1_tile_v_0_MPORT_19_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_1_tile_v_3_MPORT_19_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_1_tile_v_3_MPORT_19_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_1_tile_v_3_MPORT_19_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_1_tile_v_2_MPORT_19_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_1_tile_v_2_MPORT_19_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_1_tile_v_2_MPORT_19_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_1_tile_v_1_MPORT_19_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_1_tile_v_1_MPORT_19_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_1_tile_v_1_MPORT_19_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_1_tile_v_0_MPORT_19_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_1_tile_v_0_MPORT_19_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_1_tile_v_0_MPORT_19_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_1_MPORT_44_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_1_MPORT_44_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_1_MPORT_44_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_0_MPORT_44_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_0_MPORT_44_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_0_MPORT_44_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_1_tile_v_3_MPORT_20_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_1_tile_v_3_MPORT_20_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_1_tile_v_3_MPORT_20_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_1_tile_v_2_MPORT_20_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_1_tile_v_2_MPORT_20_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_1_tile_v_2_MPORT_20_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_1_tile_v_1_MPORT_20_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_1_tile_v_1_MPORT_20_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_1_tile_v_1_MPORT_20_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_1_tile_v_0_MPORT_20_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_1_tile_v_0_MPORT_20_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_1_tile_v_0_MPORT_20_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_1_tile_v_3_MPORT_20_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_1_tile_v_3_MPORT_20_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_1_tile_v_3_MPORT_20_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_1_tile_v_2_MPORT_20_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_1_tile_v_2_MPORT_20_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_1_tile_v_2_MPORT_20_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_1_tile_v_1_MPORT_20_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_1_tile_v_1_MPORT_20_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_1_tile_v_1_MPORT_20_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_1_tile_v_0_MPORT_20_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_1_tile_v_0_MPORT_20_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_1_tile_v_0_MPORT_20_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_3_MPORT_15_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_3_MPORT_15_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_3_MPORT_15_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_2_MPORT_15_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_2_MPORT_15_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_2_MPORT_15_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_1_MPORT_45_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_1_MPORT_45_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_1_MPORT_45_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_0_MPORT_45_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_0_MPORT_45_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_0_MPORT_45_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_1_tile_v_3_MPORT_21_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_1_tile_v_3_MPORT_21_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_1_tile_v_3_MPORT_21_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_1_tile_v_2_MPORT_21_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_1_tile_v_2_MPORT_21_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_1_tile_v_2_MPORT_21_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_1_tile_v_1_MPORT_21_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_1_tile_v_1_MPORT_21_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_1_tile_v_1_MPORT_21_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_1_tile_v_0_MPORT_21_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_1_tile_v_0_MPORT_21_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_1_tile_v_0_MPORT_21_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_1_tile_v_3_MPORT_21_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_1_tile_v_3_MPORT_21_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_1_tile_v_3_MPORT_21_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_1_tile_v_2_MPORT_21_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_1_tile_v_2_MPORT_21_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_1_tile_v_2_MPORT_21_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_1_tile_v_1_MPORT_21_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_1_tile_v_1_MPORT_21_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_1_tile_v_1_MPORT_21_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_1_tile_v_0_MPORT_21_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_1_tile_v_0_MPORT_21_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_1_tile_v_0_MPORT_21_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_1_MPORT_46_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_1_MPORT_46_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_1_MPORT_46_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_0_MPORT_46_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_0_MPORT_46_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_0_MPORT_46_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_1_tile_v_3_MPORT_22_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_1_tile_v_3_MPORT_22_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_1_tile_v_3_MPORT_22_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_1_tile_v_2_MPORT_22_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_1_tile_v_2_MPORT_22_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_1_tile_v_2_MPORT_22_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_1_tile_v_1_MPORT_22_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_1_tile_v_1_MPORT_22_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_1_tile_v_1_MPORT_22_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_1_tile_v_0_MPORT_22_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_1_tile_v_0_MPORT_22_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_1_tile_v_0_MPORT_22_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_1_tile_v_3_MPORT_22_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_1_tile_v_3_MPORT_22_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_1_tile_v_3_MPORT_22_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_1_tile_v_2_MPORT_22_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_1_tile_v_2_MPORT_22_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_1_tile_v_2_MPORT_22_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_1_tile_v_1_MPORT_22_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_1_tile_v_1_MPORT_22_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_1_tile_v_1_MPORT_22_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_1_tile_v_0_MPORT_22_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_1_tile_v_0_MPORT_22_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_1_tile_v_0_MPORT_22_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_1_MPORT_47_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_1_MPORT_47_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_1_MPORT_47_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_0_MPORT_47_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_0_MPORT_47_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_0_MPORT_47_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_1_tile_v_3_MPORT_23_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_1_tile_v_3_MPORT_23_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_1_tile_v_3_MPORT_23_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_1_tile_v_2_MPORT_23_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_1_tile_v_2_MPORT_23_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_1_tile_v_2_MPORT_23_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_1_tile_v_1_MPORT_23_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_1_tile_v_1_MPORT_23_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_1_tile_v_1_MPORT_23_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_1_tile_v_0_MPORT_23_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_1_tile_v_0_MPORT_23_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_1_tile_v_0_MPORT_23_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_1_tile_v_3_MPORT_23_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_1_tile_v_3_MPORT_23_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_1_tile_v_3_MPORT_23_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_1_tile_v_2_MPORT_23_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_1_tile_v_2_MPORT_23_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_1_tile_v_2_MPORT_23_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_1_tile_v_1_MPORT_23_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_1_tile_v_1_MPORT_23_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_1_tile_v_1_MPORT_23_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_1_tile_v_0_MPORT_23_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_1_tile_v_0_MPORT_23_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_1_tile_v_0_MPORT_23_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_1_MPORT_48_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_1_MPORT_48_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_1_MPORT_48_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_0_MPORT_48_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_0_MPORT_48_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_0_MPORT_48_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_2_tile_v_3_MPORT_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_2_tile_v_3_MPORT_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_2_tile_v_3_MPORT_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_2_tile_v_2_MPORT_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_2_tile_v_2_MPORT_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_2_tile_v_2_MPORT_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_2_tile_v_1_MPORT_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_2_tile_v_1_MPORT_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_2_tile_v_1_MPORT_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_2_tile_v_0_MPORT_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_2_tile_v_0_MPORT_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_2_tile_v_0_MPORT_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_2_tile_v_3_MPORT_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_2_tile_v_3_MPORT_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_2_tile_v_3_MPORT_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_2_tile_v_2_MPORT_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_2_tile_v_2_MPORT_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_2_tile_v_2_MPORT_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_2_tile_v_1_MPORT_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_2_tile_v_1_MPORT_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_2_tile_v_1_MPORT_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_2_tile_v_0_MPORT_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_2_tile_v_0_MPORT_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_2_tile_v_0_MPORT_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_3_MPORT_16_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_3_MPORT_16_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_3_MPORT_16_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_2_MPORT_16_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_2_MPORT_16_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_2_MPORT_16_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_1_MPORT_49_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_1_MPORT_49_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_1_MPORT_49_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_0_MPORT_49_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_0_MPORT_49_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_0_MPORT_49_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_2_tile_v_3_MPORT_1_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_2_tile_v_3_MPORT_1_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_2_tile_v_3_MPORT_1_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_2_tile_v_2_MPORT_1_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_2_tile_v_2_MPORT_1_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_2_tile_v_2_MPORT_1_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_2_tile_v_1_MPORT_1_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_2_tile_v_1_MPORT_1_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_2_tile_v_1_MPORT_1_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_2_tile_v_0_MPORT_1_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_2_tile_v_0_MPORT_1_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_2_tile_v_0_MPORT_1_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_2_tile_v_3_MPORT_1_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_2_tile_v_3_MPORT_1_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_2_tile_v_3_MPORT_1_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_2_tile_v_2_MPORT_1_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_2_tile_v_2_MPORT_1_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_2_tile_v_2_MPORT_1_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_2_tile_v_1_MPORT_1_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_2_tile_v_1_MPORT_1_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_2_tile_v_1_MPORT_1_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_2_tile_v_0_MPORT_1_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_2_tile_v_0_MPORT_1_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_2_tile_v_0_MPORT_1_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_1_MPORT_50_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_1_MPORT_50_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_1_MPORT_50_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_0_MPORT_50_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_0_MPORT_50_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_0_MPORT_50_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_2_tile_v_3_MPORT_2_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_2_tile_v_3_MPORT_2_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_2_tile_v_3_MPORT_2_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_2_tile_v_2_MPORT_2_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_2_tile_v_2_MPORT_2_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_2_tile_v_2_MPORT_2_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_2_tile_v_1_MPORT_2_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_2_tile_v_1_MPORT_2_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_2_tile_v_1_MPORT_2_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_2_tile_v_0_MPORT_2_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_2_tile_v_0_MPORT_2_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_2_tile_v_0_MPORT_2_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_2_tile_v_3_MPORT_2_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_2_tile_v_3_MPORT_2_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_2_tile_v_3_MPORT_2_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_2_tile_v_2_MPORT_2_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_2_tile_v_2_MPORT_2_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_2_tile_v_2_MPORT_2_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_2_tile_v_1_MPORT_2_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_2_tile_v_1_MPORT_2_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_2_tile_v_1_MPORT_2_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_2_tile_v_0_MPORT_2_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_2_tile_v_0_MPORT_2_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_2_tile_v_0_MPORT_2_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_3_MPORT_17_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_3_MPORT_17_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_3_MPORT_17_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_2_MPORT_17_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_2_MPORT_17_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_2_MPORT_17_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_1_MPORT_51_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_1_MPORT_51_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_1_MPORT_51_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_0_MPORT_51_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_0_MPORT_51_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_0_MPORT_51_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_2_tile_v_3_MPORT_3_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_2_tile_v_3_MPORT_3_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_2_tile_v_3_MPORT_3_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_2_tile_v_2_MPORT_3_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_2_tile_v_2_MPORT_3_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_2_tile_v_2_MPORT_3_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_2_tile_v_1_MPORT_3_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_2_tile_v_1_MPORT_3_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_2_tile_v_1_MPORT_3_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_2_tile_v_0_MPORT_3_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_2_tile_v_0_MPORT_3_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_2_tile_v_0_MPORT_3_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_2_tile_v_3_MPORT_3_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_2_tile_v_3_MPORT_3_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_2_tile_v_3_MPORT_3_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_2_tile_v_2_MPORT_3_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_2_tile_v_2_MPORT_3_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_2_tile_v_2_MPORT_3_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_2_tile_v_1_MPORT_3_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_2_tile_v_1_MPORT_3_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_2_tile_v_1_MPORT_3_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_2_tile_v_0_MPORT_3_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_2_tile_v_0_MPORT_3_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_2_tile_v_0_MPORT_3_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_1_MPORT_52_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_1_MPORT_52_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_1_MPORT_52_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_0_MPORT_52_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_0_MPORT_52_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_0_MPORT_52_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_2_tile_v_3_MPORT_4_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_2_tile_v_3_MPORT_4_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_2_tile_v_3_MPORT_4_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_2_tile_v_2_MPORT_4_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_2_tile_v_2_MPORT_4_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_2_tile_v_2_MPORT_4_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_2_tile_v_1_MPORT_4_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_2_tile_v_1_MPORT_4_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_2_tile_v_1_MPORT_4_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_2_tile_v_0_MPORT_4_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_2_tile_v_0_MPORT_4_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_2_tile_v_0_MPORT_4_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_2_tile_v_3_MPORT_4_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_2_tile_v_3_MPORT_4_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_2_tile_v_3_MPORT_4_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_2_tile_v_2_MPORT_4_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_2_tile_v_2_MPORT_4_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_2_tile_v_2_MPORT_4_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_2_tile_v_1_MPORT_4_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_2_tile_v_1_MPORT_4_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_2_tile_v_1_MPORT_4_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_2_tile_v_0_MPORT_4_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_2_tile_v_0_MPORT_4_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_2_tile_v_0_MPORT_4_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_1_MPORT_53_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_1_MPORT_53_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_1_MPORT_53_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_0_MPORT_53_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_0_MPORT_53_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_0_MPORT_53_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_2_tile_v_3_MPORT_5_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_2_tile_v_3_MPORT_5_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_2_tile_v_3_MPORT_5_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_2_tile_v_2_MPORT_5_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_2_tile_v_2_MPORT_5_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_2_tile_v_2_MPORT_5_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_2_tile_v_1_MPORT_5_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_2_tile_v_1_MPORT_5_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_2_tile_v_1_MPORT_5_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_2_tile_v_0_MPORT_5_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_2_tile_v_0_MPORT_5_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_2_tile_v_0_MPORT_5_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_2_tile_v_3_MPORT_5_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_2_tile_v_3_MPORT_5_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_2_tile_v_3_MPORT_5_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_2_tile_v_2_MPORT_5_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_2_tile_v_2_MPORT_5_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_2_tile_v_2_MPORT_5_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_2_tile_v_1_MPORT_5_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_2_tile_v_1_MPORT_5_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_2_tile_v_1_MPORT_5_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_2_tile_v_0_MPORT_5_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_2_tile_v_0_MPORT_5_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_2_tile_v_0_MPORT_5_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_1_MPORT_54_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_1_MPORT_54_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_1_MPORT_54_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_0_MPORT_54_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_0_MPORT_54_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_0_MPORT_54_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_2_tile_v_3_MPORT_6_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_2_tile_v_3_MPORT_6_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_2_tile_v_3_MPORT_6_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_2_tile_v_2_MPORT_6_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_2_tile_v_2_MPORT_6_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_2_tile_v_2_MPORT_6_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_2_tile_v_1_MPORT_6_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_2_tile_v_1_MPORT_6_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_2_tile_v_1_MPORT_6_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_2_tile_v_0_MPORT_6_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_2_tile_v_0_MPORT_6_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_2_tile_v_0_MPORT_6_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_2_tile_v_3_MPORT_6_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_2_tile_v_3_MPORT_6_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_2_tile_v_3_MPORT_6_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_2_tile_v_2_MPORT_6_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_2_tile_v_2_MPORT_6_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_2_tile_v_2_MPORT_6_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_2_tile_v_1_MPORT_6_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_2_tile_v_1_MPORT_6_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_2_tile_v_1_MPORT_6_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_2_tile_v_0_MPORT_6_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_2_tile_v_0_MPORT_6_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_2_tile_v_0_MPORT_6_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_3_MPORT_18_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_3_MPORT_18_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_3_MPORT_18_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_2_MPORT_18_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_2_MPORT_18_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_2_MPORT_18_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_1_MPORT_55_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_1_MPORT_55_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_1_MPORT_55_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_0_MPORT_55_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_0_MPORT_55_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_0_MPORT_55_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_2_tile_v_3_MPORT_7_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_2_tile_v_3_MPORT_7_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_2_tile_v_3_MPORT_7_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_2_tile_v_2_MPORT_7_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_2_tile_v_2_MPORT_7_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_2_tile_v_2_MPORT_7_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_2_tile_v_1_MPORT_7_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_2_tile_v_1_MPORT_7_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_2_tile_v_1_MPORT_7_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_2_tile_v_0_MPORT_7_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_2_tile_v_0_MPORT_7_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_2_tile_v_0_MPORT_7_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_2_tile_v_3_MPORT_7_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_2_tile_v_3_MPORT_7_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_2_tile_v_3_MPORT_7_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_2_tile_v_2_MPORT_7_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_2_tile_v_2_MPORT_7_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_2_tile_v_2_MPORT_7_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_2_tile_v_1_MPORT_7_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_2_tile_v_1_MPORT_7_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_2_tile_v_1_MPORT_7_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_2_tile_v_0_MPORT_7_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_2_tile_v_0_MPORT_7_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_2_tile_v_0_MPORT_7_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_1_MPORT_56_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_1_MPORT_56_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_1_MPORT_56_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_0_MPORT_56_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_0_MPORT_56_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_0_MPORT_56_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_2_tile_v_3_MPORT_8_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_2_tile_v_3_MPORT_8_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_2_tile_v_3_MPORT_8_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_2_tile_v_2_MPORT_8_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_2_tile_v_2_MPORT_8_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_2_tile_v_2_MPORT_8_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_2_tile_v_1_MPORT_8_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_2_tile_v_1_MPORT_8_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_2_tile_v_1_MPORT_8_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_2_tile_v_0_MPORT_8_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_2_tile_v_0_MPORT_8_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_2_tile_v_0_MPORT_8_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_2_tile_v_3_MPORT_8_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_2_tile_v_3_MPORT_8_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_2_tile_v_3_MPORT_8_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_2_tile_v_2_MPORT_8_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_2_tile_v_2_MPORT_8_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_2_tile_v_2_MPORT_8_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_2_tile_v_1_MPORT_8_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_2_tile_v_1_MPORT_8_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_2_tile_v_1_MPORT_8_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_2_tile_v_0_MPORT_8_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_2_tile_v_0_MPORT_8_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_2_tile_v_0_MPORT_8_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_3_MPORT_19_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_3_MPORT_19_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_3_MPORT_19_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_2_MPORT_19_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_2_MPORT_19_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_2_MPORT_19_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_1_MPORT_57_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_1_MPORT_57_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_1_MPORT_57_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_0_MPORT_57_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_0_MPORT_57_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_0_MPORT_57_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_2_tile_v_3_MPORT_9_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_2_tile_v_3_MPORT_9_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_2_tile_v_3_MPORT_9_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_2_tile_v_2_MPORT_9_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_2_tile_v_2_MPORT_9_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_2_tile_v_2_MPORT_9_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_2_tile_v_1_MPORT_9_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_2_tile_v_1_MPORT_9_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_2_tile_v_1_MPORT_9_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_2_tile_v_0_MPORT_9_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_2_tile_v_0_MPORT_9_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_2_tile_v_0_MPORT_9_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_2_tile_v_3_MPORT_9_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_2_tile_v_3_MPORT_9_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_2_tile_v_3_MPORT_9_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_2_tile_v_2_MPORT_9_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_2_tile_v_2_MPORT_9_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_2_tile_v_2_MPORT_9_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_2_tile_v_1_MPORT_9_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_2_tile_v_1_MPORT_9_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_2_tile_v_1_MPORT_9_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_2_tile_v_0_MPORT_9_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_2_tile_v_0_MPORT_9_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_2_tile_v_0_MPORT_9_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_1_MPORT_58_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_1_MPORT_58_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_1_MPORT_58_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_0_MPORT_58_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_0_MPORT_58_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_0_MPORT_58_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_2_tile_v_3_MPORT_10_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_2_tile_v_3_MPORT_10_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_2_tile_v_3_MPORT_10_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_2_tile_v_2_MPORT_10_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_2_tile_v_2_MPORT_10_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_2_tile_v_2_MPORT_10_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_2_tile_v_1_MPORT_10_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_2_tile_v_1_MPORT_10_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_2_tile_v_1_MPORT_10_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_2_tile_v_0_MPORT_10_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_2_tile_v_0_MPORT_10_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_2_tile_v_0_MPORT_10_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_2_tile_v_3_MPORT_10_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_2_tile_v_3_MPORT_10_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_2_tile_v_3_MPORT_10_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_2_tile_v_2_MPORT_10_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_2_tile_v_2_MPORT_10_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_2_tile_v_2_MPORT_10_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_2_tile_v_1_MPORT_10_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_2_tile_v_1_MPORT_10_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_2_tile_v_1_MPORT_10_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_2_tile_v_0_MPORT_10_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_2_tile_v_0_MPORT_10_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_2_tile_v_0_MPORT_10_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_1_MPORT_59_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_1_MPORT_59_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_1_MPORT_59_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_0_MPORT_59_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_0_MPORT_59_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_0_MPORT_59_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_2_tile_v_3_MPORT_11_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_2_tile_v_3_MPORT_11_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_2_tile_v_3_MPORT_11_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_2_tile_v_2_MPORT_11_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_2_tile_v_2_MPORT_11_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_2_tile_v_2_MPORT_11_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_2_tile_v_1_MPORT_11_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_2_tile_v_1_MPORT_11_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_2_tile_v_1_MPORT_11_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_2_tile_v_0_MPORT_11_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_2_tile_v_0_MPORT_11_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_2_tile_v_0_MPORT_11_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_2_tile_v_3_MPORT_11_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_2_tile_v_3_MPORT_11_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_2_tile_v_3_MPORT_11_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_2_tile_v_2_MPORT_11_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_2_tile_v_2_MPORT_11_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_2_tile_v_2_MPORT_11_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_2_tile_v_1_MPORT_11_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_2_tile_v_1_MPORT_11_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_2_tile_v_1_MPORT_11_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_2_tile_v_0_MPORT_11_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_2_tile_v_0_MPORT_11_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_2_tile_v_0_MPORT_11_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_1_MPORT_60_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_1_MPORT_60_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_1_MPORT_60_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_0_MPORT_60_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_0_MPORT_60_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_0_MPORT_60_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_2_tile_v_3_MPORT_12_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_2_tile_v_3_MPORT_12_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_2_tile_v_3_MPORT_12_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_2_tile_v_2_MPORT_12_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_2_tile_v_2_MPORT_12_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_2_tile_v_2_MPORT_12_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_2_tile_v_1_MPORT_12_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_2_tile_v_1_MPORT_12_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_2_tile_v_1_MPORT_12_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_2_tile_v_0_MPORT_12_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_2_tile_v_0_MPORT_12_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_2_tile_v_0_MPORT_12_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_2_tile_v_3_MPORT_12_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_2_tile_v_3_MPORT_12_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_2_tile_v_3_MPORT_12_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_2_tile_v_2_MPORT_12_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_2_tile_v_2_MPORT_12_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_2_tile_v_2_MPORT_12_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_2_tile_v_1_MPORT_12_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_2_tile_v_1_MPORT_12_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_2_tile_v_1_MPORT_12_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_2_tile_v_0_MPORT_12_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_2_tile_v_0_MPORT_12_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_2_tile_v_0_MPORT_12_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_3_MPORT_20_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_3_MPORT_20_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_3_MPORT_20_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_2_MPORT_20_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_2_MPORT_20_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_2_MPORT_20_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_1_MPORT_61_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_1_MPORT_61_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_1_MPORT_61_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_0_MPORT_61_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_0_MPORT_61_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_0_MPORT_61_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_2_tile_v_3_MPORT_13_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_2_tile_v_3_MPORT_13_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_2_tile_v_3_MPORT_13_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_2_tile_v_2_MPORT_13_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_2_tile_v_2_MPORT_13_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_2_tile_v_2_MPORT_13_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_2_tile_v_1_MPORT_13_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_2_tile_v_1_MPORT_13_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_2_tile_v_1_MPORT_13_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_2_tile_v_0_MPORT_13_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_2_tile_v_0_MPORT_13_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_2_tile_v_0_MPORT_13_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_2_tile_v_3_MPORT_13_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_2_tile_v_3_MPORT_13_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_2_tile_v_3_MPORT_13_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_2_tile_v_2_MPORT_13_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_2_tile_v_2_MPORT_13_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_2_tile_v_2_MPORT_13_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_2_tile_v_1_MPORT_13_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_2_tile_v_1_MPORT_13_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_2_tile_v_1_MPORT_13_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_2_tile_v_0_MPORT_13_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_2_tile_v_0_MPORT_13_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_2_tile_v_0_MPORT_13_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_1_MPORT_62_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_1_MPORT_62_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_1_MPORT_62_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_0_MPORT_62_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_0_MPORT_62_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_0_MPORT_62_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_2_tile_v_3_MPORT_14_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_2_tile_v_3_MPORT_14_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_2_tile_v_3_MPORT_14_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_2_tile_v_2_MPORT_14_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_2_tile_v_2_MPORT_14_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_2_tile_v_2_MPORT_14_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_2_tile_v_1_MPORT_14_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_2_tile_v_1_MPORT_14_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_2_tile_v_1_MPORT_14_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_2_tile_v_0_MPORT_14_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_2_tile_v_0_MPORT_14_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_2_tile_v_0_MPORT_14_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_2_tile_v_3_MPORT_14_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_2_tile_v_3_MPORT_14_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_2_tile_v_3_MPORT_14_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_2_tile_v_2_MPORT_14_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_2_tile_v_2_MPORT_14_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_2_tile_v_2_MPORT_14_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_2_tile_v_1_MPORT_14_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_2_tile_v_1_MPORT_14_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_2_tile_v_1_MPORT_14_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_2_tile_v_0_MPORT_14_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_2_tile_v_0_MPORT_14_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_2_tile_v_0_MPORT_14_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_3_MPORT_21_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_3_MPORT_21_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_3_MPORT_21_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_2_MPORT_21_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_2_MPORT_21_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_2_MPORT_21_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_1_MPORT_63_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_1_MPORT_63_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_1_MPORT_63_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_0_MPORT_63_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_0_MPORT_63_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_0_MPORT_63_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_2_tile_v_3_MPORT_15_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_2_tile_v_3_MPORT_15_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_2_tile_v_3_MPORT_15_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_2_tile_v_2_MPORT_15_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_2_tile_v_2_MPORT_15_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_2_tile_v_2_MPORT_15_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_2_tile_v_1_MPORT_15_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_2_tile_v_1_MPORT_15_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_2_tile_v_1_MPORT_15_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_2_tile_v_0_MPORT_15_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_2_tile_v_0_MPORT_15_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_2_tile_v_0_MPORT_15_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_2_tile_v_3_MPORT_15_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_2_tile_v_3_MPORT_15_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_2_tile_v_3_MPORT_15_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_2_tile_v_2_MPORT_15_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_2_tile_v_2_MPORT_15_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_2_tile_v_2_MPORT_15_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_2_tile_v_1_MPORT_15_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_2_tile_v_1_MPORT_15_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_2_tile_v_1_MPORT_15_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_2_tile_v_0_MPORT_15_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_2_tile_v_0_MPORT_15_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_2_tile_v_0_MPORT_15_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_1_MPORT_64_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_1_MPORT_64_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_1_MPORT_64_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_0_MPORT_64_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_0_MPORT_64_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_0_MPORT_64_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_2_tile_v_3_MPORT_16_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_2_tile_v_3_MPORT_16_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_2_tile_v_3_MPORT_16_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_2_tile_v_2_MPORT_16_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_2_tile_v_2_MPORT_16_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_2_tile_v_2_MPORT_16_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_2_tile_v_1_MPORT_16_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_2_tile_v_1_MPORT_16_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_2_tile_v_1_MPORT_16_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_2_tile_v_0_MPORT_16_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_2_tile_v_0_MPORT_16_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_2_tile_v_0_MPORT_16_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_2_tile_v_3_MPORT_16_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_2_tile_v_3_MPORT_16_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_2_tile_v_3_MPORT_16_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_2_tile_v_2_MPORT_16_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_2_tile_v_2_MPORT_16_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_2_tile_v_2_MPORT_16_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_2_tile_v_1_MPORT_16_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_2_tile_v_1_MPORT_16_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_2_tile_v_1_MPORT_16_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_2_tile_v_0_MPORT_16_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_2_tile_v_0_MPORT_16_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_2_tile_v_0_MPORT_16_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_1_MPORT_65_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_1_MPORT_65_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_1_MPORT_65_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_0_MPORT_65_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_0_MPORT_65_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_0_MPORT_65_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_2_tile_v_3_MPORT_17_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_2_tile_v_3_MPORT_17_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_2_tile_v_3_MPORT_17_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_2_tile_v_2_MPORT_17_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_2_tile_v_2_MPORT_17_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_2_tile_v_2_MPORT_17_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_2_tile_v_1_MPORT_17_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_2_tile_v_1_MPORT_17_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_2_tile_v_1_MPORT_17_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_2_tile_v_0_MPORT_17_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_2_tile_v_0_MPORT_17_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_2_tile_v_0_MPORT_17_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_2_tile_v_3_MPORT_17_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_2_tile_v_3_MPORT_17_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_2_tile_v_3_MPORT_17_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_2_tile_v_2_MPORT_17_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_2_tile_v_2_MPORT_17_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_2_tile_v_2_MPORT_17_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_2_tile_v_1_MPORT_17_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_2_tile_v_1_MPORT_17_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_2_tile_v_1_MPORT_17_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_2_tile_v_0_MPORT_17_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_2_tile_v_0_MPORT_17_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_2_tile_v_0_MPORT_17_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_1_MPORT_66_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_1_MPORT_66_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_1_MPORT_66_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_0_MPORT_66_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_0_MPORT_66_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_0_MPORT_66_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_2_tile_v_3_MPORT_18_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_2_tile_v_3_MPORT_18_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_2_tile_v_3_MPORT_18_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_2_tile_v_2_MPORT_18_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_2_tile_v_2_MPORT_18_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_2_tile_v_2_MPORT_18_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_2_tile_v_1_MPORT_18_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_2_tile_v_1_MPORT_18_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_2_tile_v_1_MPORT_18_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_2_tile_v_0_MPORT_18_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_2_tile_v_0_MPORT_18_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_2_tile_v_0_MPORT_18_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_2_tile_v_3_MPORT_18_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_2_tile_v_3_MPORT_18_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_2_tile_v_3_MPORT_18_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_2_tile_v_2_MPORT_18_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_2_tile_v_2_MPORT_18_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_2_tile_v_2_MPORT_18_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_2_tile_v_1_MPORT_18_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_2_tile_v_1_MPORT_18_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_2_tile_v_1_MPORT_18_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_2_tile_v_0_MPORT_18_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_2_tile_v_0_MPORT_18_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_2_tile_v_0_MPORT_18_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_3_MPORT_22_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_3_MPORT_22_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_3_MPORT_22_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_2_MPORT_22_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_2_MPORT_22_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_2_MPORT_22_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_1_MPORT_67_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_1_MPORT_67_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_1_MPORT_67_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_0_MPORT_67_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_0_MPORT_67_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_0_MPORT_67_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_2_tile_v_3_MPORT_19_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_2_tile_v_3_MPORT_19_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_2_tile_v_3_MPORT_19_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_2_tile_v_2_MPORT_19_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_2_tile_v_2_MPORT_19_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_2_tile_v_2_MPORT_19_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_2_tile_v_1_MPORT_19_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_2_tile_v_1_MPORT_19_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_2_tile_v_1_MPORT_19_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_2_tile_v_0_MPORT_19_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_2_tile_v_0_MPORT_19_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_2_tile_v_0_MPORT_19_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_2_tile_v_3_MPORT_19_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_2_tile_v_3_MPORT_19_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_2_tile_v_3_MPORT_19_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_2_tile_v_2_MPORT_19_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_2_tile_v_2_MPORT_19_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_2_tile_v_2_MPORT_19_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_2_tile_v_1_MPORT_19_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_2_tile_v_1_MPORT_19_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_2_tile_v_1_MPORT_19_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_2_tile_v_0_MPORT_19_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_2_tile_v_0_MPORT_19_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_2_tile_v_0_MPORT_19_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_1_MPORT_68_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_1_MPORT_68_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_1_MPORT_68_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_0_MPORT_68_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_0_MPORT_68_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_0_MPORT_68_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_2_tile_v_3_MPORT_20_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_2_tile_v_3_MPORT_20_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_2_tile_v_3_MPORT_20_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_2_tile_v_2_MPORT_20_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_2_tile_v_2_MPORT_20_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_2_tile_v_2_MPORT_20_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_2_tile_v_1_MPORT_20_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_2_tile_v_1_MPORT_20_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_2_tile_v_1_MPORT_20_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_2_tile_v_0_MPORT_20_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_2_tile_v_0_MPORT_20_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_2_tile_v_0_MPORT_20_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_2_tile_v_3_MPORT_20_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_2_tile_v_3_MPORT_20_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_2_tile_v_3_MPORT_20_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_2_tile_v_2_MPORT_20_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_2_tile_v_2_MPORT_20_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_2_tile_v_2_MPORT_20_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_2_tile_v_1_MPORT_20_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_2_tile_v_1_MPORT_20_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_2_tile_v_1_MPORT_20_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_2_tile_v_0_MPORT_20_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_2_tile_v_0_MPORT_20_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_2_tile_v_0_MPORT_20_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_3_MPORT_23_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_3_MPORT_23_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_3_MPORT_23_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_2_MPORT_23_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_2_MPORT_23_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_2_MPORT_23_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_1_MPORT_69_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_1_MPORT_69_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_1_MPORT_69_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_0_MPORT_69_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_0_MPORT_69_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_0_MPORT_69_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_2_tile_v_3_MPORT_21_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_2_tile_v_3_MPORT_21_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_2_tile_v_3_MPORT_21_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_2_tile_v_2_MPORT_21_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_2_tile_v_2_MPORT_21_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_2_tile_v_2_MPORT_21_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_2_tile_v_1_MPORT_21_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_2_tile_v_1_MPORT_21_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_2_tile_v_1_MPORT_21_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_2_tile_v_0_MPORT_21_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_2_tile_v_0_MPORT_21_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_2_tile_v_0_MPORT_21_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_2_tile_v_3_MPORT_21_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_2_tile_v_3_MPORT_21_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_2_tile_v_3_MPORT_21_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_2_tile_v_2_MPORT_21_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_2_tile_v_2_MPORT_21_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_2_tile_v_2_MPORT_21_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_2_tile_v_1_MPORT_21_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_2_tile_v_1_MPORT_21_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_2_tile_v_1_MPORT_21_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_2_tile_v_0_MPORT_21_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_2_tile_v_0_MPORT_21_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_2_tile_v_0_MPORT_21_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_1_MPORT_70_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_1_MPORT_70_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_1_MPORT_70_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_0_MPORT_70_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_0_MPORT_70_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_0_MPORT_70_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_2_tile_v_3_MPORT_22_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_2_tile_v_3_MPORT_22_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_2_tile_v_3_MPORT_22_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_2_tile_v_2_MPORT_22_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_2_tile_v_2_MPORT_22_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_2_tile_v_2_MPORT_22_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_2_tile_v_1_MPORT_22_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_2_tile_v_1_MPORT_22_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_2_tile_v_1_MPORT_22_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_2_tile_v_0_MPORT_22_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_2_tile_v_0_MPORT_22_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_2_tile_v_0_MPORT_22_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_2_tile_v_3_MPORT_22_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_2_tile_v_3_MPORT_22_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_2_tile_v_3_MPORT_22_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_2_tile_v_2_MPORT_22_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_2_tile_v_2_MPORT_22_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_2_tile_v_2_MPORT_22_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_2_tile_v_1_MPORT_22_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_2_tile_v_1_MPORT_22_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_2_tile_v_1_MPORT_22_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_2_tile_v_0_MPORT_22_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_2_tile_v_0_MPORT_22_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_2_tile_v_0_MPORT_22_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_1_MPORT_71_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_1_MPORT_71_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_1_MPORT_71_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_0_MPORT_71_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_0_MPORT_71_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_0_MPORT_71_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_2_tile_v_3_MPORT_23_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_2_tile_v_3_MPORT_23_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_2_tile_v_3_MPORT_23_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_2_tile_v_2_MPORT_23_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_2_tile_v_2_MPORT_23_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_2_tile_v_2_MPORT_23_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_2_tile_v_1_MPORT_23_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_2_tile_v_1_MPORT_23_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_2_tile_v_1_MPORT_23_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_2_tile_v_0_MPORT_23_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_2_tile_v_0_MPORT_23_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_2_tile_v_0_MPORT_23_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_2_tile_v_3_MPORT_23_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_2_tile_v_3_MPORT_23_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_2_tile_v_3_MPORT_23_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_2_tile_v_2_MPORT_23_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_2_tile_v_2_MPORT_23_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_2_tile_v_2_MPORT_23_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_2_tile_v_1_MPORT_23_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_2_tile_v_1_MPORT_23_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_2_tile_v_1_MPORT_23_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_2_tile_v_0_MPORT_23_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_2_tile_v_0_MPORT_23_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_2_tile_v_0_MPORT_23_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_1_MPORT_72_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_1_MPORT_72_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_1_MPORT_72_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_0_MPORT_72_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_0_MPORT_72_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_0_MPORT_72_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_3_tile_v_3_MPORT_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_3_tile_v_3_MPORT_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_3_tile_v_3_MPORT_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_3_tile_v_2_MPORT_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_3_tile_v_2_MPORT_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_3_tile_v_2_MPORT_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_3_tile_v_1_MPORT_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_3_tile_v_1_MPORT_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_3_tile_v_1_MPORT_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_3_tile_v_0_MPORT_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_3_tile_v_0_MPORT_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_3_tile_v_0_MPORT_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_3_tile_v_3_MPORT_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_3_tile_v_3_MPORT_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_3_tile_v_3_MPORT_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_3_tile_v_2_MPORT_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_3_tile_v_2_MPORT_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_3_tile_v_2_MPORT_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_3_tile_v_1_MPORT_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_3_tile_v_1_MPORT_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_3_tile_v_1_MPORT_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_3_tile_v_0_MPORT_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_3_tile_v_0_MPORT_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_3_tile_v_0_MPORT_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_3_MPORT_24_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_3_MPORT_24_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_3_MPORT_24_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_2_MPORT_24_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_2_MPORT_24_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_2_MPORT_24_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_1_MPORT_73_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_1_MPORT_73_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_1_MPORT_73_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_0_MPORT_73_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_0_MPORT_73_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_0_MPORT_73_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_3_tile_v_3_MPORT_1_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_3_tile_v_3_MPORT_1_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_3_tile_v_3_MPORT_1_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_3_tile_v_2_MPORT_1_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_3_tile_v_2_MPORT_1_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_3_tile_v_2_MPORT_1_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_3_tile_v_1_MPORT_1_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_3_tile_v_1_MPORT_1_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_3_tile_v_1_MPORT_1_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_3_tile_v_0_MPORT_1_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_3_tile_v_0_MPORT_1_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_3_tile_v_0_MPORT_1_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_3_tile_v_3_MPORT_1_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_3_tile_v_3_MPORT_1_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_3_tile_v_3_MPORT_1_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_3_tile_v_2_MPORT_1_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_3_tile_v_2_MPORT_1_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_3_tile_v_2_MPORT_1_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_3_tile_v_1_MPORT_1_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_3_tile_v_1_MPORT_1_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_3_tile_v_1_MPORT_1_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_3_tile_v_0_MPORT_1_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_3_tile_v_0_MPORT_1_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_3_tile_v_0_MPORT_1_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_1_MPORT_74_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_1_MPORT_74_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_1_MPORT_74_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_0_MPORT_74_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_0_MPORT_74_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_0_MPORT_74_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_3_tile_v_3_MPORT_2_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_3_tile_v_3_MPORT_2_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_3_tile_v_3_MPORT_2_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_3_tile_v_2_MPORT_2_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_3_tile_v_2_MPORT_2_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_3_tile_v_2_MPORT_2_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_3_tile_v_1_MPORT_2_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_3_tile_v_1_MPORT_2_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_3_tile_v_1_MPORT_2_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_3_tile_v_0_MPORT_2_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_3_tile_v_0_MPORT_2_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_3_tile_v_0_MPORT_2_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_3_tile_v_3_MPORT_2_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_3_tile_v_3_MPORT_2_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_3_tile_v_3_MPORT_2_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_3_tile_v_2_MPORT_2_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_3_tile_v_2_MPORT_2_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_3_tile_v_2_MPORT_2_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_3_tile_v_1_MPORT_2_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_3_tile_v_1_MPORT_2_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_3_tile_v_1_MPORT_2_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_3_tile_v_0_MPORT_2_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_3_tile_v_0_MPORT_2_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_3_tile_v_0_MPORT_2_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_3_MPORT_25_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_3_MPORT_25_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_3_MPORT_25_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_2_MPORT_25_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_2_MPORT_25_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_2_MPORT_25_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_1_MPORT_75_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_1_MPORT_75_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_1_MPORT_75_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_0_MPORT_75_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_0_MPORT_75_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_0_MPORT_75_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_3_tile_v_3_MPORT_3_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_3_tile_v_3_MPORT_3_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_3_tile_v_3_MPORT_3_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_3_tile_v_2_MPORT_3_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_3_tile_v_2_MPORT_3_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_3_tile_v_2_MPORT_3_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_3_tile_v_1_MPORT_3_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_3_tile_v_1_MPORT_3_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_3_tile_v_1_MPORT_3_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_3_tile_v_0_MPORT_3_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_3_tile_v_0_MPORT_3_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_3_tile_v_0_MPORT_3_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_3_tile_v_3_MPORT_3_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_3_tile_v_3_MPORT_3_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_3_tile_v_3_MPORT_3_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_3_tile_v_2_MPORT_3_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_3_tile_v_2_MPORT_3_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_3_tile_v_2_MPORT_3_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_3_tile_v_1_MPORT_3_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_3_tile_v_1_MPORT_3_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_3_tile_v_1_MPORT_3_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_3_tile_v_0_MPORT_3_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_3_tile_v_0_MPORT_3_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_3_tile_v_0_MPORT_3_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_1_MPORT_76_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_1_MPORT_76_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_1_MPORT_76_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_0_MPORT_76_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_0_MPORT_76_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_0_MPORT_76_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_3_tile_v_3_MPORT_4_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_3_tile_v_3_MPORT_4_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_3_tile_v_3_MPORT_4_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_3_tile_v_2_MPORT_4_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_3_tile_v_2_MPORT_4_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_3_tile_v_2_MPORT_4_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_3_tile_v_1_MPORT_4_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_3_tile_v_1_MPORT_4_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_3_tile_v_1_MPORT_4_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_3_tile_v_0_MPORT_4_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_3_tile_v_0_MPORT_4_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_3_tile_v_0_MPORT_4_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_3_tile_v_3_MPORT_4_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_3_tile_v_3_MPORT_4_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_3_tile_v_3_MPORT_4_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_3_tile_v_2_MPORT_4_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_3_tile_v_2_MPORT_4_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_3_tile_v_2_MPORT_4_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_3_tile_v_1_MPORT_4_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_3_tile_v_1_MPORT_4_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_3_tile_v_1_MPORT_4_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_3_tile_v_0_MPORT_4_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_3_tile_v_0_MPORT_4_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_3_tile_v_0_MPORT_4_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_1_MPORT_77_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_1_MPORT_77_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_1_MPORT_77_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_0_MPORT_77_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_0_MPORT_77_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_0_MPORT_77_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_3_tile_v_3_MPORT_5_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_3_tile_v_3_MPORT_5_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_3_tile_v_3_MPORT_5_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_3_tile_v_2_MPORT_5_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_3_tile_v_2_MPORT_5_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_3_tile_v_2_MPORT_5_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_3_tile_v_1_MPORT_5_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_3_tile_v_1_MPORT_5_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_3_tile_v_1_MPORT_5_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_3_tile_v_0_MPORT_5_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_3_tile_v_0_MPORT_5_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_3_tile_v_0_MPORT_5_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_3_tile_v_3_MPORT_5_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_3_tile_v_3_MPORT_5_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_3_tile_v_3_MPORT_5_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_3_tile_v_2_MPORT_5_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_3_tile_v_2_MPORT_5_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_3_tile_v_2_MPORT_5_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_3_tile_v_1_MPORT_5_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_3_tile_v_1_MPORT_5_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_3_tile_v_1_MPORT_5_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_3_tile_v_0_MPORT_5_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_3_tile_v_0_MPORT_5_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_3_tile_v_0_MPORT_5_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_1_MPORT_78_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_1_MPORT_78_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_1_MPORT_78_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_0_MPORT_78_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_0_MPORT_78_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_0_MPORT_78_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_3_tile_v_3_MPORT_6_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_3_tile_v_3_MPORT_6_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_3_tile_v_3_MPORT_6_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_3_tile_v_2_MPORT_6_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_3_tile_v_2_MPORT_6_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_3_tile_v_2_MPORT_6_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_3_tile_v_1_MPORT_6_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_3_tile_v_1_MPORT_6_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_3_tile_v_1_MPORT_6_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_3_tile_v_0_MPORT_6_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_3_tile_v_0_MPORT_6_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_3_tile_v_0_MPORT_6_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_3_tile_v_3_MPORT_6_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_3_tile_v_3_MPORT_6_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_3_tile_v_3_MPORT_6_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_3_tile_v_2_MPORT_6_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_3_tile_v_2_MPORT_6_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_3_tile_v_2_MPORT_6_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_3_tile_v_1_MPORT_6_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_3_tile_v_1_MPORT_6_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_3_tile_v_1_MPORT_6_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_3_tile_v_0_MPORT_6_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_3_tile_v_0_MPORT_6_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_3_tile_v_0_MPORT_6_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_3_MPORT_26_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_3_MPORT_26_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_3_MPORT_26_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_2_MPORT_26_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_2_MPORT_26_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_2_MPORT_26_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_1_MPORT_79_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_1_MPORT_79_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_1_MPORT_79_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_0_MPORT_79_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_0_MPORT_79_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_0_MPORT_79_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_3_tile_v_3_MPORT_7_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_3_tile_v_3_MPORT_7_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_3_tile_v_3_MPORT_7_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_3_tile_v_2_MPORT_7_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_3_tile_v_2_MPORT_7_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_3_tile_v_2_MPORT_7_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_3_tile_v_1_MPORT_7_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_3_tile_v_1_MPORT_7_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_3_tile_v_1_MPORT_7_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_3_tile_v_0_MPORT_7_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_3_tile_v_0_MPORT_7_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_3_tile_v_0_MPORT_7_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_3_tile_v_3_MPORT_7_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_3_tile_v_3_MPORT_7_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_3_tile_v_3_MPORT_7_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_3_tile_v_2_MPORT_7_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_3_tile_v_2_MPORT_7_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_3_tile_v_2_MPORT_7_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_3_tile_v_1_MPORT_7_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_3_tile_v_1_MPORT_7_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_3_tile_v_1_MPORT_7_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_3_tile_v_0_MPORT_7_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_3_tile_v_0_MPORT_7_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_3_tile_v_0_MPORT_7_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_1_MPORT_80_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_1_MPORT_80_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_1_MPORT_80_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_0_MPORT_80_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_0_MPORT_80_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_0_MPORT_80_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_3_tile_v_3_MPORT_8_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_3_tile_v_3_MPORT_8_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_3_tile_v_3_MPORT_8_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_3_tile_v_2_MPORT_8_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_3_tile_v_2_MPORT_8_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_3_tile_v_2_MPORT_8_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_3_tile_v_1_MPORT_8_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_3_tile_v_1_MPORT_8_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_3_tile_v_1_MPORT_8_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_3_tile_v_0_MPORT_8_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_3_tile_v_0_MPORT_8_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_3_tile_v_0_MPORT_8_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_3_tile_v_3_MPORT_8_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_3_tile_v_3_MPORT_8_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_3_tile_v_3_MPORT_8_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_3_tile_v_2_MPORT_8_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_3_tile_v_2_MPORT_8_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_3_tile_v_2_MPORT_8_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_3_tile_v_1_MPORT_8_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_3_tile_v_1_MPORT_8_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_3_tile_v_1_MPORT_8_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_3_tile_v_0_MPORT_8_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_3_tile_v_0_MPORT_8_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_3_tile_v_0_MPORT_8_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_3_MPORT_27_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_3_MPORT_27_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_3_MPORT_27_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_2_MPORT_27_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_2_MPORT_27_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_2_MPORT_27_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_1_MPORT_81_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_1_MPORT_81_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_1_MPORT_81_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_0_MPORT_81_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_0_MPORT_81_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_0_MPORT_81_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_3_tile_v_3_MPORT_9_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_3_tile_v_3_MPORT_9_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_3_tile_v_3_MPORT_9_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_3_tile_v_2_MPORT_9_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_3_tile_v_2_MPORT_9_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_3_tile_v_2_MPORT_9_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_3_tile_v_1_MPORT_9_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_3_tile_v_1_MPORT_9_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_3_tile_v_1_MPORT_9_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_3_tile_v_0_MPORT_9_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_3_tile_v_0_MPORT_9_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_3_tile_v_0_MPORT_9_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_3_tile_v_3_MPORT_9_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_3_tile_v_3_MPORT_9_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_3_tile_v_3_MPORT_9_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_3_tile_v_2_MPORT_9_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_3_tile_v_2_MPORT_9_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_3_tile_v_2_MPORT_9_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_3_tile_v_1_MPORT_9_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_3_tile_v_1_MPORT_9_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_3_tile_v_1_MPORT_9_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_3_tile_v_0_MPORT_9_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_3_tile_v_0_MPORT_9_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_3_tile_v_0_MPORT_9_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_1_MPORT_82_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_1_MPORT_82_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_1_MPORT_82_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_0_MPORT_82_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_0_MPORT_82_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_0_MPORT_82_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_3_tile_v_3_MPORT_10_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_3_tile_v_3_MPORT_10_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_3_tile_v_3_MPORT_10_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_3_tile_v_2_MPORT_10_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_3_tile_v_2_MPORT_10_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_3_tile_v_2_MPORT_10_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_3_tile_v_1_MPORT_10_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_3_tile_v_1_MPORT_10_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_3_tile_v_1_MPORT_10_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_3_tile_v_0_MPORT_10_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_3_tile_v_0_MPORT_10_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_3_tile_v_0_MPORT_10_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_3_tile_v_3_MPORT_10_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_3_tile_v_3_MPORT_10_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_3_tile_v_3_MPORT_10_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_3_tile_v_2_MPORT_10_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_3_tile_v_2_MPORT_10_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_3_tile_v_2_MPORT_10_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_3_tile_v_1_MPORT_10_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_3_tile_v_1_MPORT_10_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_3_tile_v_1_MPORT_10_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_3_tile_v_0_MPORT_10_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_3_tile_v_0_MPORT_10_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_3_tile_v_0_MPORT_10_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_1_MPORT_83_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_1_MPORT_83_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_1_MPORT_83_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_0_MPORT_83_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_0_MPORT_83_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_0_MPORT_83_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_3_tile_v_3_MPORT_11_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_3_tile_v_3_MPORT_11_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_3_tile_v_3_MPORT_11_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_3_tile_v_2_MPORT_11_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_3_tile_v_2_MPORT_11_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_3_tile_v_2_MPORT_11_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_3_tile_v_1_MPORT_11_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_3_tile_v_1_MPORT_11_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_3_tile_v_1_MPORT_11_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_3_tile_v_0_MPORT_11_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_3_tile_v_0_MPORT_11_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_3_tile_v_0_MPORT_11_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_3_tile_v_3_MPORT_11_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_3_tile_v_3_MPORT_11_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_3_tile_v_3_MPORT_11_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_3_tile_v_2_MPORT_11_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_3_tile_v_2_MPORT_11_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_3_tile_v_2_MPORT_11_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_3_tile_v_1_MPORT_11_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_3_tile_v_1_MPORT_11_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_3_tile_v_1_MPORT_11_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_3_tile_v_0_MPORT_11_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_3_tile_v_0_MPORT_11_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_3_tile_v_0_MPORT_11_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_1_MPORT_84_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_1_MPORT_84_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_1_MPORT_84_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_0_MPORT_84_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_0_MPORT_84_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_0_MPORT_84_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_3_tile_v_3_MPORT_12_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_3_tile_v_3_MPORT_12_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_3_tile_v_3_MPORT_12_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_3_tile_v_2_MPORT_12_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_3_tile_v_2_MPORT_12_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_3_tile_v_2_MPORT_12_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_3_tile_v_1_MPORT_12_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_3_tile_v_1_MPORT_12_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_3_tile_v_1_MPORT_12_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_3_tile_v_0_MPORT_12_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_3_tile_v_0_MPORT_12_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_3_tile_v_0_MPORT_12_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_3_tile_v_3_MPORT_12_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_3_tile_v_3_MPORT_12_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_3_tile_v_3_MPORT_12_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_3_tile_v_2_MPORT_12_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_3_tile_v_2_MPORT_12_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_3_tile_v_2_MPORT_12_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_3_tile_v_1_MPORT_12_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_3_tile_v_1_MPORT_12_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_3_tile_v_1_MPORT_12_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_3_tile_v_0_MPORT_12_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_3_tile_v_0_MPORT_12_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_3_tile_v_0_MPORT_12_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_3_MPORT_28_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_3_MPORT_28_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_3_MPORT_28_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_2_MPORT_28_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_2_MPORT_28_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_2_MPORT_28_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_1_MPORT_85_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_1_MPORT_85_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_1_MPORT_85_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_0_MPORT_85_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_0_MPORT_85_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_0_MPORT_85_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_3_tile_v_3_MPORT_13_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_3_tile_v_3_MPORT_13_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_3_tile_v_3_MPORT_13_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_3_tile_v_2_MPORT_13_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_3_tile_v_2_MPORT_13_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_3_tile_v_2_MPORT_13_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_3_tile_v_1_MPORT_13_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_3_tile_v_1_MPORT_13_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_3_tile_v_1_MPORT_13_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_3_tile_v_0_MPORT_13_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_3_tile_v_0_MPORT_13_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_3_tile_v_0_MPORT_13_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_3_tile_v_3_MPORT_13_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_3_tile_v_3_MPORT_13_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_3_tile_v_3_MPORT_13_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_3_tile_v_2_MPORT_13_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_3_tile_v_2_MPORT_13_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_3_tile_v_2_MPORT_13_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_3_tile_v_1_MPORT_13_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_3_tile_v_1_MPORT_13_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_3_tile_v_1_MPORT_13_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_3_tile_v_0_MPORT_13_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_3_tile_v_0_MPORT_13_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_3_tile_v_0_MPORT_13_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_1_MPORT_86_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_1_MPORT_86_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_1_MPORT_86_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_0_MPORT_86_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_0_MPORT_86_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_0_MPORT_86_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_3_tile_v_3_MPORT_14_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_3_tile_v_3_MPORT_14_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_3_tile_v_3_MPORT_14_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_3_tile_v_2_MPORT_14_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_3_tile_v_2_MPORT_14_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_3_tile_v_2_MPORT_14_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_3_tile_v_1_MPORT_14_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_3_tile_v_1_MPORT_14_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_3_tile_v_1_MPORT_14_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_3_tile_v_0_MPORT_14_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_3_tile_v_0_MPORT_14_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_3_tile_v_0_MPORT_14_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_3_tile_v_3_MPORT_14_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_3_tile_v_3_MPORT_14_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_3_tile_v_3_MPORT_14_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_3_tile_v_2_MPORT_14_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_3_tile_v_2_MPORT_14_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_3_tile_v_2_MPORT_14_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_3_tile_v_1_MPORT_14_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_3_tile_v_1_MPORT_14_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_3_tile_v_1_MPORT_14_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_3_tile_v_0_MPORT_14_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_3_tile_v_0_MPORT_14_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_3_tile_v_0_MPORT_14_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_3_MPORT_29_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_3_MPORT_29_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_3_MPORT_29_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_2_MPORT_29_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_2_MPORT_29_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_2_MPORT_29_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_1_MPORT_87_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_1_MPORT_87_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_1_MPORT_87_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_0_MPORT_87_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_0_MPORT_87_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_0_MPORT_87_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_3_tile_v_3_MPORT_15_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_3_tile_v_3_MPORT_15_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_3_tile_v_3_MPORT_15_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_3_tile_v_2_MPORT_15_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_3_tile_v_2_MPORT_15_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_3_tile_v_2_MPORT_15_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_3_tile_v_1_MPORT_15_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_3_tile_v_1_MPORT_15_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_3_tile_v_1_MPORT_15_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_3_tile_v_0_MPORT_15_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_3_tile_v_0_MPORT_15_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_3_tile_v_0_MPORT_15_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_3_tile_v_3_MPORT_15_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_3_tile_v_3_MPORT_15_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_3_tile_v_3_MPORT_15_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_3_tile_v_2_MPORT_15_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_3_tile_v_2_MPORT_15_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_3_tile_v_2_MPORT_15_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_3_tile_v_1_MPORT_15_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_3_tile_v_1_MPORT_15_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_3_tile_v_1_MPORT_15_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_3_tile_v_0_MPORT_15_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_3_tile_v_0_MPORT_15_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_3_tile_v_0_MPORT_15_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_1_MPORT_88_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_1_MPORT_88_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_1_MPORT_88_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_0_MPORT_88_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_0_MPORT_88_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_0_MPORT_88_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_3_tile_v_3_MPORT_16_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_3_tile_v_3_MPORT_16_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_3_tile_v_3_MPORT_16_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_3_tile_v_2_MPORT_16_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_3_tile_v_2_MPORT_16_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_3_tile_v_2_MPORT_16_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_3_tile_v_1_MPORT_16_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_3_tile_v_1_MPORT_16_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_3_tile_v_1_MPORT_16_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_3_tile_v_0_MPORT_16_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_3_tile_v_0_MPORT_16_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_3_tile_v_0_MPORT_16_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_3_tile_v_3_MPORT_16_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_3_tile_v_3_MPORT_16_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_3_tile_v_3_MPORT_16_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_3_tile_v_2_MPORT_16_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_3_tile_v_2_MPORT_16_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_3_tile_v_2_MPORT_16_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_3_tile_v_1_MPORT_16_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_3_tile_v_1_MPORT_16_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_3_tile_v_1_MPORT_16_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_3_tile_v_0_MPORT_16_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_3_tile_v_0_MPORT_16_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_3_tile_v_0_MPORT_16_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_1_MPORT_89_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_1_MPORT_89_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_1_MPORT_89_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_0_MPORT_89_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_0_MPORT_89_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_0_MPORT_89_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_3_tile_v_3_MPORT_17_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_3_tile_v_3_MPORT_17_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_3_tile_v_3_MPORT_17_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_3_tile_v_2_MPORT_17_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_3_tile_v_2_MPORT_17_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_3_tile_v_2_MPORT_17_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_3_tile_v_1_MPORT_17_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_3_tile_v_1_MPORT_17_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_3_tile_v_1_MPORT_17_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_3_tile_v_0_MPORT_17_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_3_tile_v_0_MPORT_17_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_3_tile_v_0_MPORT_17_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_3_tile_v_3_MPORT_17_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_3_tile_v_3_MPORT_17_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_3_tile_v_3_MPORT_17_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_3_tile_v_2_MPORT_17_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_3_tile_v_2_MPORT_17_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_3_tile_v_2_MPORT_17_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_3_tile_v_1_MPORT_17_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_3_tile_v_1_MPORT_17_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_3_tile_v_1_MPORT_17_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_3_tile_v_0_MPORT_17_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_3_tile_v_0_MPORT_17_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_3_tile_v_0_MPORT_17_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_1_MPORT_90_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_1_MPORT_90_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_1_MPORT_90_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_0_MPORT_90_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_0_MPORT_90_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_0_MPORT_90_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_3_tile_v_3_MPORT_18_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_3_tile_v_3_MPORT_18_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_3_tile_v_3_MPORT_18_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_3_tile_v_2_MPORT_18_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_3_tile_v_2_MPORT_18_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_3_tile_v_2_MPORT_18_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_3_tile_v_1_MPORT_18_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_3_tile_v_1_MPORT_18_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_3_tile_v_1_MPORT_18_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_3_tile_v_0_MPORT_18_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_3_tile_v_0_MPORT_18_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_3_tile_v_0_MPORT_18_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_3_tile_v_3_MPORT_18_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_3_tile_v_3_MPORT_18_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_3_tile_v_3_MPORT_18_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_3_tile_v_2_MPORT_18_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_3_tile_v_2_MPORT_18_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_3_tile_v_2_MPORT_18_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_3_tile_v_1_MPORT_18_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_3_tile_v_1_MPORT_18_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_3_tile_v_1_MPORT_18_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_3_tile_v_0_MPORT_18_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_3_tile_v_0_MPORT_18_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_3_tile_v_0_MPORT_18_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_3_MPORT_30_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_3_MPORT_30_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_3_MPORT_30_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_2_MPORT_30_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_2_MPORT_30_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_2_MPORT_30_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_1_MPORT_91_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_1_MPORT_91_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_1_MPORT_91_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_0_MPORT_91_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_0_MPORT_91_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_0_MPORT_91_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_3_tile_v_3_MPORT_19_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_3_tile_v_3_MPORT_19_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_3_tile_v_3_MPORT_19_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_3_tile_v_2_MPORT_19_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_3_tile_v_2_MPORT_19_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_3_tile_v_2_MPORT_19_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_3_tile_v_1_MPORT_19_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_3_tile_v_1_MPORT_19_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_3_tile_v_1_MPORT_19_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_3_tile_v_0_MPORT_19_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_3_tile_v_0_MPORT_19_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_3_tile_v_0_MPORT_19_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_3_tile_v_3_MPORT_19_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_3_tile_v_3_MPORT_19_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_3_tile_v_3_MPORT_19_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_3_tile_v_2_MPORT_19_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_3_tile_v_2_MPORT_19_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_3_tile_v_2_MPORT_19_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_3_tile_v_1_MPORT_19_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_3_tile_v_1_MPORT_19_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_3_tile_v_1_MPORT_19_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_3_tile_v_0_MPORT_19_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_3_tile_v_0_MPORT_19_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_3_tile_v_0_MPORT_19_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_1_MPORT_92_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_1_MPORT_92_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_1_MPORT_92_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_0_MPORT_92_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_0_MPORT_92_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_0_MPORT_92_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_3_tile_v_3_MPORT_20_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_3_tile_v_3_MPORT_20_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_3_tile_v_3_MPORT_20_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_3_tile_v_2_MPORT_20_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_3_tile_v_2_MPORT_20_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_3_tile_v_2_MPORT_20_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_3_tile_v_1_MPORT_20_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_3_tile_v_1_MPORT_20_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_3_tile_v_1_MPORT_20_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_3_tile_v_0_MPORT_20_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_3_tile_v_0_MPORT_20_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_3_tile_v_0_MPORT_20_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_3_tile_v_3_MPORT_20_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_3_tile_v_3_MPORT_20_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_3_tile_v_3_MPORT_20_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_3_tile_v_2_MPORT_20_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_3_tile_v_2_MPORT_20_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_3_tile_v_2_MPORT_20_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_3_tile_v_1_MPORT_20_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_3_tile_v_1_MPORT_20_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_3_tile_v_1_MPORT_20_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_3_tile_v_0_MPORT_20_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_3_tile_v_0_MPORT_20_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_3_tile_v_0_MPORT_20_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_3_MPORT_31_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_3_MPORT_31_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_3_MPORT_31_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_2_MPORT_31_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_2_MPORT_31_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_2_MPORT_31_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_1_MPORT_93_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_1_MPORT_93_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_1_MPORT_93_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_0_MPORT_93_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_0_MPORT_93_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_0_MPORT_93_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_3_tile_v_3_MPORT_21_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_3_tile_v_3_MPORT_21_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_3_tile_v_3_MPORT_21_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_3_tile_v_2_MPORT_21_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_3_tile_v_2_MPORT_21_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_3_tile_v_2_MPORT_21_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_3_tile_v_1_MPORT_21_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_3_tile_v_1_MPORT_21_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_3_tile_v_1_MPORT_21_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_3_tile_v_0_MPORT_21_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_3_tile_v_0_MPORT_21_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_3_tile_v_0_MPORT_21_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_3_tile_v_3_MPORT_21_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_3_tile_v_3_MPORT_21_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_3_tile_v_3_MPORT_21_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_3_tile_v_2_MPORT_21_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_3_tile_v_2_MPORT_21_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_3_tile_v_2_MPORT_21_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_3_tile_v_1_MPORT_21_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_3_tile_v_1_MPORT_21_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_3_tile_v_1_MPORT_21_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_3_tile_v_0_MPORT_21_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_3_tile_v_0_MPORT_21_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_3_tile_v_0_MPORT_21_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_1_MPORT_94_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_1_MPORT_94_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_1_MPORT_94_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_0_MPORT_94_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_0_MPORT_94_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_0_MPORT_94_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_3_tile_v_3_MPORT_22_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_3_tile_v_3_MPORT_22_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_3_tile_v_3_MPORT_22_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_3_tile_v_2_MPORT_22_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_3_tile_v_2_MPORT_22_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_3_tile_v_2_MPORT_22_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_3_tile_v_1_MPORT_22_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_3_tile_v_1_MPORT_22_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_3_tile_v_1_MPORT_22_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_3_tile_v_0_MPORT_22_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_3_tile_v_0_MPORT_22_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_3_tile_v_0_MPORT_22_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_3_tile_v_3_MPORT_22_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_3_tile_v_3_MPORT_22_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_3_tile_v_3_MPORT_22_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_3_tile_v_2_MPORT_22_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_3_tile_v_2_MPORT_22_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_3_tile_v_2_MPORT_22_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_3_tile_v_1_MPORT_22_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_3_tile_v_1_MPORT_22_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_3_tile_v_1_MPORT_22_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_3_tile_v_0_MPORT_22_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_3_tile_v_0_MPORT_22_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_3_tile_v_0_MPORT_22_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_1_MPORT_95_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_1_MPORT_95_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_1_MPORT_95_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_0_MPORT_95_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_0_MPORT_95_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_0_MPORT_95_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_3_tile_v_3_MPORT_23_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_3_tile_v_3_MPORT_23_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_3_tile_v_3_MPORT_23_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_3_tile_v_2_MPORT_23_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_3_tile_v_2_MPORT_23_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_3_tile_v_2_MPORT_23_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_3_tile_v_1_MPORT_23_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_3_tile_v_1_MPORT_23_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_3_tile_v_1_MPORT_23_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_3_tile_v_0_MPORT_23_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_3_tile_v_0_MPORT_23_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_3_tile_v_0_MPORT_23_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_3_tile_v_3_MPORT_23_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_3_tile_v_3_MPORT_23_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_3_tile_v_3_MPORT_23_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_3_tile_v_2_MPORT_23_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_3_tile_v_2_MPORT_23_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_3_tile_v_2_MPORT_23_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_3_tile_v_1_MPORT_23_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_3_tile_v_1_MPORT_23_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_3_tile_v_1_MPORT_23_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_3_tile_v_0_MPORT_23_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_3_tile_v_0_MPORT_23_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_3_tile_v_0_MPORT_23_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_1_MPORT_96_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_1_MPORT_96_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_1_MPORT_96_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_0_MPORT_96_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_0_MPORT_96_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_0_MPORT_96_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_4_tile_v_3_MPORT_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_4_tile_v_3_MPORT_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_4_tile_v_3_MPORT_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_4_tile_v_2_MPORT_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_4_tile_v_2_MPORT_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_4_tile_v_2_MPORT_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_4_tile_v_1_MPORT_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_4_tile_v_1_MPORT_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_4_tile_v_1_MPORT_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_4_tile_v_0_MPORT_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_4_tile_v_0_MPORT_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_4_tile_v_0_MPORT_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_4_tile_v_3_MPORT_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_4_tile_v_3_MPORT_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_4_tile_v_3_MPORT_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_4_tile_v_2_MPORT_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_4_tile_v_2_MPORT_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_4_tile_v_2_MPORT_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_4_tile_v_1_MPORT_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_4_tile_v_1_MPORT_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_4_tile_v_1_MPORT_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_4_tile_v_0_MPORT_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_4_tile_v_0_MPORT_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_4_tile_v_0_MPORT_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_3_MPORT_32_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_3_MPORT_32_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_3_MPORT_32_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_2_MPORT_32_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_2_MPORT_32_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_2_MPORT_32_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_1_MPORT_97_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_1_MPORT_97_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_1_MPORT_97_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_0_MPORT_97_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_0_MPORT_97_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_0_MPORT_97_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_4_tile_v_3_MPORT_1_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_4_tile_v_3_MPORT_1_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_4_tile_v_3_MPORT_1_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_4_tile_v_2_MPORT_1_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_4_tile_v_2_MPORT_1_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_4_tile_v_2_MPORT_1_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_4_tile_v_1_MPORT_1_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_4_tile_v_1_MPORT_1_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_4_tile_v_1_MPORT_1_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_4_tile_v_0_MPORT_1_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_4_tile_v_0_MPORT_1_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_4_tile_v_0_MPORT_1_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_4_tile_v_3_MPORT_1_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_4_tile_v_3_MPORT_1_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_4_tile_v_3_MPORT_1_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_4_tile_v_2_MPORT_1_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_4_tile_v_2_MPORT_1_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_4_tile_v_2_MPORT_1_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_4_tile_v_1_MPORT_1_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_4_tile_v_1_MPORT_1_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_4_tile_v_1_MPORT_1_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_4_tile_v_0_MPORT_1_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_4_tile_v_0_MPORT_1_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_4_tile_v_0_MPORT_1_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_1_MPORT_98_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_1_MPORT_98_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_1_MPORT_98_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_0_MPORT_98_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_0_MPORT_98_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_0_MPORT_98_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_4_tile_v_3_MPORT_2_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_4_tile_v_3_MPORT_2_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_4_tile_v_3_MPORT_2_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_4_tile_v_2_MPORT_2_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_4_tile_v_2_MPORT_2_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_4_tile_v_2_MPORT_2_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_4_tile_v_1_MPORT_2_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_4_tile_v_1_MPORT_2_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_4_tile_v_1_MPORT_2_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_4_tile_v_0_MPORT_2_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_4_tile_v_0_MPORT_2_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_4_tile_v_0_MPORT_2_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_4_tile_v_3_MPORT_2_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_4_tile_v_3_MPORT_2_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_4_tile_v_3_MPORT_2_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_4_tile_v_2_MPORT_2_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_4_tile_v_2_MPORT_2_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_4_tile_v_2_MPORT_2_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_4_tile_v_1_MPORT_2_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_4_tile_v_1_MPORT_2_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_4_tile_v_1_MPORT_2_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_4_tile_v_0_MPORT_2_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_4_tile_v_0_MPORT_2_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_4_tile_v_0_MPORT_2_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_3_MPORT_33_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_3_MPORT_33_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_3_MPORT_33_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_2_MPORT_33_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_2_MPORT_33_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_2_MPORT_33_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_1_MPORT_99_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_1_MPORT_99_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_1_MPORT_99_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_0_MPORT_99_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_0_MPORT_99_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_0_MPORT_99_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_4_tile_v_3_MPORT_3_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_4_tile_v_3_MPORT_3_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_4_tile_v_3_MPORT_3_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_4_tile_v_2_MPORT_3_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_4_tile_v_2_MPORT_3_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_4_tile_v_2_MPORT_3_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_4_tile_v_1_MPORT_3_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_4_tile_v_1_MPORT_3_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_4_tile_v_1_MPORT_3_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_4_tile_v_0_MPORT_3_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_4_tile_v_0_MPORT_3_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_4_tile_v_0_MPORT_3_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_4_tile_v_3_MPORT_3_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_4_tile_v_3_MPORT_3_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_4_tile_v_3_MPORT_3_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_4_tile_v_2_MPORT_3_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_4_tile_v_2_MPORT_3_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_4_tile_v_2_MPORT_3_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_4_tile_v_1_MPORT_3_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_4_tile_v_1_MPORT_3_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_4_tile_v_1_MPORT_3_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_4_tile_v_0_MPORT_3_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_4_tile_v_0_MPORT_3_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_4_tile_v_0_MPORT_3_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_1_MPORT_100_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_1_MPORT_100_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_1_MPORT_100_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_0_MPORT_100_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_0_MPORT_100_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_0_MPORT_100_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_4_tile_v_3_MPORT_4_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_4_tile_v_3_MPORT_4_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_4_tile_v_3_MPORT_4_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_4_tile_v_2_MPORT_4_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_4_tile_v_2_MPORT_4_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_4_tile_v_2_MPORT_4_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_4_tile_v_1_MPORT_4_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_4_tile_v_1_MPORT_4_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_4_tile_v_1_MPORT_4_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_4_tile_v_0_MPORT_4_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_4_tile_v_0_MPORT_4_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_4_tile_v_0_MPORT_4_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_4_tile_v_3_MPORT_4_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_4_tile_v_3_MPORT_4_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_4_tile_v_3_MPORT_4_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_4_tile_v_2_MPORT_4_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_4_tile_v_2_MPORT_4_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_4_tile_v_2_MPORT_4_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_4_tile_v_1_MPORT_4_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_4_tile_v_1_MPORT_4_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_4_tile_v_1_MPORT_4_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_4_tile_v_0_MPORT_4_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_4_tile_v_0_MPORT_4_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_4_tile_v_0_MPORT_4_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_1_MPORT_101_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_1_MPORT_101_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_1_MPORT_101_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_0_MPORT_101_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_0_MPORT_101_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_0_MPORT_101_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_4_tile_v_3_MPORT_5_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_4_tile_v_3_MPORT_5_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_4_tile_v_3_MPORT_5_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_4_tile_v_2_MPORT_5_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_4_tile_v_2_MPORT_5_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_4_tile_v_2_MPORT_5_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_4_tile_v_1_MPORT_5_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_4_tile_v_1_MPORT_5_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_4_tile_v_1_MPORT_5_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_4_tile_v_0_MPORT_5_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_4_tile_v_0_MPORT_5_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_4_tile_v_0_MPORT_5_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_4_tile_v_3_MPORT_5_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_4_tile_v_3_MPORT_5_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_4_tile_v_3_MPORT_5_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_4_tile_v_2_MPORT_5_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_4_tile_v_2_MPORT_5_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_4_tile_v_2_MPORT_5_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_4_tile_v_1_MPORT_5_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_4_tile_v_1_MPORT_5_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_4_tile_v_1_MPORT_5_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_4_tile_v_0_MPORT_5_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_4_tile_v_0_MPORT_5_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_4_tile_v_0_MPORT_5_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_1_MPORT_102_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_1_MPORT_102_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_1_MPORT_102_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_0_MPORT_102_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_0_MPORT_102_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_0_MPORT_102_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_4_tile_v_3_MPORT_6_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_4_tile_v_3_MPORT_6_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_4_tile_v_3_MPORT_6_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_4_tile_v_2_MPORT_6_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_4_tile_v_2_MPORT_6_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_4_tile_v_2_MPORT_6_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_4_tile_v_1_MPORT_6_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_4_tile_v_1_MPORT_6_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_4_tile_v_1_MPORT_6_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_4_tile_v_0_MPORT_6_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_4_tile_v_0_MPORT_6_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_4_tile_v_0_MPORT_6_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_4_tile_v_3_MPORT_6_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_4_tile_v_3_MPORT_6_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_4_tile_v_3_MPORT_6_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_4_tile_v_2_MPORT_6_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_4_tile_v_2_MPORT_6_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_4_tile_v_2_MPORT_6_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_4_tile_v_1_MPORT_6_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_4_tile_v_1_MPORT_6_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_4_tile_v_1_MPORT_6_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_4_tile_v_0_MPORT_6_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_4_tile_v_0_MPORT_6_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_4_tile_v_0_MPORT_6_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_3_MPORT_34_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_3_MPORT_34_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_3_MPORT_34_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_2_MPORT_34_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_2_MPORT_34_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_2_MPORT_34_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_1_MPORT_103_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_1_MPORT_103_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_1_MPORT_103_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_0_MPORT_103_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_0_MPORT_103_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_0_MPORT_103_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_4_tile_v_3_MPORT_7_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_4_tile_v_3_MPORT_7_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_4_tile_v_3_MPORT_7_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_4_tile_v_2_MPORT_7_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_4_tile_v_2_MPORT_7_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_4_tile_v_2_MPORT_7_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_4_tile_v_1_MPORT_7_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_4_tile_v_1_MPORT_7_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_4_tile_v_1_MPORT_7_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_4_tile_v_0_MPORT_7_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_4_tile_v_0_MPORT_7_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_4_tile_v_0_MPORT_7_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_4_tile_v_3_MPORT_7_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_4_tile_v_3_MPORT_7_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_4_tile_v_3_MPORT_7_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_4_tile_v_2_MPORT_7_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_4_tile_v_2_MPORT_7_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_4_tile_v_2_MPORT_7_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_4_tile_v_1_MPORT_7_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_4_tile_v_1_MPORT_7_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_4_tile_v_1_MPORT_7_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_4_tile_v_0_MPORT_7_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_4_tile_v_0_MPORT_7_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_4_tile_v_0_MPORT_7_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_1_MPORT_104_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_1_MPORT_104_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_1_MPORT_104_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_0_MPORT_104_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_0_MPORT_104_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_0_MPORT_104_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_4_tile_v_3_MPORT_8_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_4_tile_v_3_MPORT_8_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_4_tile_v_3_MPORT_8_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_4_tile_v_2_MPORT_8_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_4_tile_v_2_MPORT_8_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_4_tile_v_2_MPORT_8_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_4_tile_v_1_MPORT_8_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_4_tile_v_1_MPORT_8_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_4_tile_v_1_MPORT_8_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_4_tile_v_0_MPORT_8_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_4_tile_v_0_MPORT_8_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_4_tile_v_0_MPORT_8_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_4_tile_v_3_MPORT_8_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_4_tile_v_3_MPORT_8_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_4_tile_v_3_MPORT_8_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_4_tile_v_2_MPORT_8_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_4_tile_v_2_MPORT_8_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_4_tile_v_2_MPORT_8_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_4_tile_v_1_MPORT_8_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_4_tile_v_1_MPORT_8_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_4_tile_v_1_MPORT_8_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_4_tile_v_0_MPORT_8_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_4_tile_v_0_MPORT_8_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_4_tile_v_0_MPORT_8_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_3_MPORT_35_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_3_MPORT_35_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_3_MPORT_35_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_2_MPORT_35_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_2_MPORT_35_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_2_MPORT_35_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_1_MPORT_105_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_1_MPORT_105_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_1_MPORT_105_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_0_MPORT_105_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_0_MPORT_105_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_0_MPORT_105_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_4_tile_v_3_MPORT_9_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_4_tile_v_3_MPORT_9_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_4_tile_v_3_MPORT_9_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_4_tile_v_2_MPORT_9_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_4_tile_v_2_MPORT_9_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_4_tile_v_2_MPORT_9_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_4_tile_v_1_MPORT_9_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_4_tile_v_1_MPORT_9_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_4_tile_v_1_MPORT_9_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_4_tile_v_0_MPORT_9_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_4_tile_v_0_MPORT_9_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_4_tile_v_0_MPORT_9_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_4_tile_v_3_MPORT_9_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_4_tile_v_3_MPORT_9_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_4_tile_v_3_MPORT_9_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_4_tile_v_2_MPORT_9_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_4_tile_v_2_MPORT_9_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_4_tile_v_2_MPORT_9_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_4_tile_v_1_MPORT_9_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_4_tile_v_1_MPORT_9_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_4_tile_v_1_MPORT_9_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_4_tile_v_0_MPORT_9_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_4_tile_v_0_MPORT_9_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_4_tile_v_0_MPORT_9_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_1_MPORT_106_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_1_MPORT_106_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_1_MPORT_106_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_0_MPORT_106_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_0_MPORT_106_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_0_MPORT_106_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_4_tile_v_3_MPORT_10_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_4_tile_v_3_MPORT_10_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_4_tile_v_3_MPORT_10_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_4_tile_v_2_MPORT_10_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_4_tile_v_2_MPORT_10_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_4_tile_v_2_MPORT_10_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_4_tile_v_1_MPORT_10_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_4_tile_v_1_MPORT_10_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_4_tile_v_1_MPORT_10_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_4_tile_v_0_MPORT_10_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_4_tile_v_0_MPORT_10_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_4_tile_v_0_MPORT_10_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_4_tile_v_3_MPORT_10_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_4_tile_v_3_MPORT_10_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_4_tile_v_3_MPORT_10_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_4_tile_v_2_MPORT_10_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_4_tile_v_2_MPORT_10_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_4_tile_v_2_MPORT_10_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_4_tile_v_1_MPORT_10_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_4_tile_v_1_MPORT_10_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_4_tile_v_1_MPORT_10_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_4_tile_v_0_MPORT_10_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_4_tile_v_0_MPORT_10_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_4_tile_v_0_MPORT_10_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_1_MPORT_107_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_1_MPORT_107_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_1_MPORT_107_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_0_MPORT_107_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_0_MPORT_107_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_0_MPORT_107_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_4_tile_v_3_MPORT_11_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_4_tile_v_3_MPORT_11_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_4_tile_v_3_MPORT_11_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_4_tile_v_2_MPORT_11_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_4_tile_v_2_MPORT_11_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_4_tile_v_2_MPORT_11_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_4_tile_v_1_MPORT_11_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_4_tile_v_1_MPORT_11_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_4_tile_v_1_MPORT_11_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_4_tile_v_0_MPORT_11_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_4_tile_v_0_MPORT_11_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_4_tile_v_0_MPORT_11_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_4_tile_v_3_MPORT_11_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_4_tile_v_3_MPORT_11_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_4_tile_v_3_MPORT_11_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_4_tile_v_2_MPORT_11_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_4_tile_v_2_MPORT_11_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_4_tile_v_2_MPORT_11_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_4_tile_v_1_MPORT_11_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_4_tile_v_1_MPORT_11_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_4_tile_v_1_MPORT_11_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_4_tile_v_0_MPORT_11_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_4_tile_v_0_MPORT_11_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_4_tile_v_0_MPORT_11_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_1_MPORT_108_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_1_MPORT_108_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_1_MPORT_108_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_0_MPORT_108_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_0_MPORT_108_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_0_MPORT_108_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_4_tile_v_3_MPORT_12_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_4_tile_v_3_MPORT_12_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_4_tile_v_3_MPORT_12_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_4_tile_v_2_MPORT_12_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_4_tile_v_2_MPORT_12_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_4_tile_v_2_MPORT_12_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_4_tile_v_1_MPORT_12_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_4_tile_v_1_MPORT_12_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_4_tile_v_1_MPORT_12_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_4_tile_v_0_MPORT_12_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_4_tile_v_0_MPORT_12_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_4_tile_v_0_MPORT_12_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_4_tile_v_3_MPORT_12_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_4_tile_v_3_MPORT_12_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_4_tile_v_3_MPORT_12_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_4_tile_v_2_MPORT_12_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_4_tile_v_2_MPORT_12_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_4_tile_v_2_MPORT_12_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_4_tile_v_1_MPORT_12_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_4_tile_v_1_MPORT_12_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_4_tile_v_1_MPORT_12_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_4_tile_v_0_MPORT_12_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_4_tile_v_0_MPORT_12_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_4_tile_v_0_MPORT_12_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_3_MPORT_36_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_3_MPORT_36_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_3_MPORT_36_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_2_MPORT_36_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_2_MPORT_36_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_2_MPORT_36_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_1_MPORT_109_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_1_MPORT_109_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_1_MPORT_109_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_0_MPORT_109_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_0_MPORT_109_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_0_MPORT_109_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_4_tile_v_3_MPORT_13_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_4_tile_v_3_MPORT_13_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_4_tile_v_3_MPORT_13_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_4_tile_v_2_MPORT_13_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_4_tile_v_2_MPORT_13_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_4_tile_v_2_MPORT_13_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_4_tile_v_1_MPORT_13_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_4_tile_v_1_MPORT_13_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_4_tile_v_1_MPORT_13_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_4_tile_v_0_MPORT_13_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_4_tile_v_0_MPORT_13_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_4_tile_v_0_MPORT_13_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_4_tile_v_3_MPORT_13_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_4_tile_v_3_MPORT_13_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_4_tile_v_3_MPORT_13_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_4_tile_v_2_MPORT_13_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_4_tile_v_2_MPORT_13_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_4_tile_v_2_MPORT_13_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_4_tile_v_1_MPORT_13_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_4_tile_v_1_MPORT_13_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_4_tile_v_1_MPORT_13_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_4_tile_v_0_MPORT_13_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_4_tile_v_0_MPORT_13_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_4_tile_v_0_MPORT_13_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_1_MPORT_110_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_1_MPORT_110_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_1_MPORT_110_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_0_MPORT_110_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_0_MPORT_110_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_0_MPORT_110_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_4_tile_v_3_MPORT_14_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_4_tile_v_3_MPORT_14_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_4_tile_v_3_MPORT_14_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_4_tile_v_2_MPORT_14_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_4_tile_v_2_MPORT_14_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_4_tile_v_2_MPORT_14_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_4_tile_v_1_MPORT_14_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_4_tile_v_1_MPORT_14_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_4_tile_v_1_MPORT_14_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_4_tile_v_0_MPORT_14_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_4_tile_v_0_MPORT_14_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_4_tile_v_0_MPORT_14_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_4_tile_v_3_MPORT_14_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_4_tile_v_3_MPORT_14_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_4_tile_v_3_MPORT_14_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_4_tile_v_2_MPORT_14_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_4_tile_v_2_MPORT_14_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_4_tile_v_2_MPORT_14_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_4_tile_v_1_MPORT_14_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_4_tile_v_1_MPORT_14_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_4_tile_v_1_MPORT_14_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_4_tile_v_0_MPORT_14_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_4_tile_v_0_MPORT_14_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_4_tile_v_0_MPORT_14_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_3_MPORT_37_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_3_MPORT_37_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_3_MPORT_37_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_2_MPORT_37_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_2_MPORT_37_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_2_MPORT_37_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_1_MPORT_111_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_1_MPORT_111_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_1_MPORT_111_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_0_MPORT_111_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_0_MPORT_111_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_0_MPORT_111_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_4_tile_v_3_MPORT_15_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_4_tile_v_3_MPORT_15_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_4_tile_v_3_MPORT_15_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_4_tile_v_2_MPORT_15_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_4_tile_v_2_MPORT_15_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_4_tile_v_2_MPORT_15_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_4_tile_v_1_MPORT_15_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_4_tile_v_1_MPORT_15_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_4_tile_v_1_MPORT_15_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_4_tile_v_0_MPORT_15_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_4_tile_v_0_MPORT_15_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_4_tile_v_0_MPORT_15_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_4_tile_v_3_MPORT_15_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_4_tile_v_3_MPORT_15_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_4_tile_v_3_MPORT_15_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_4_tile_v_2_MPORT_15_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_4_tile_v_2_MPORT_15_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_4_tile_v_2_MPORT_15_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_4_tile_v_1_MPORT_15_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_4_tile_v_1_MPORT_15_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_4_tile_v_1_MPORT_15_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_4_tile_v_0_MPORT_15_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_4_tile_v_0_MPORT_15_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_4_tile_v_0_MPORT_15_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_1_MPORT_112_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_1_MPORT_112_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_1_MPORT_112_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_0_MPORT_112_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_0_MPORT_112_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_0_MPORT_112_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_4_tile_v_3_MPORT_16_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_4_tile_v_3_MPORT_16_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_4_tile_v_3_MPORT_16_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_4_tile_v_2_MPORT_16_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_4_tile_v_2_MPORT_16_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_4_tile_v_2_MPORT_16_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_4_tile_v_1_MPORT_16_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_4_tile_v_1_MPORT_16_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_4_tile_v_1_MPORT_16_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_4_tile_v_0_MPORT_16_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_4_tile_v_0_MPORT_16_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_4_tile_v_0_MPORT_16_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_4_tile_v_3_MPORT_16_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_4_tile_v_3_MPORT_16_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_4_tile_v_3_MPORT_16_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_4_tile_v_2_MPORT_16_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_4_tile_v_2_MPORT_16_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_4_tile_v_2_MPORT_16_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_4_tile_v_1_MPORT_16_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_4_tile_v_1_MPORT_16_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_4_tile_v_1_MPORT_16_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_4_tile_v_0_MPORT_16_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_4_tile_v_0_MPORT_16_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_4_tile_v_0_MPORT_16_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_1_MPORT_113_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_1_MPORT_113_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_1_MPORT_113_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_0_MPORT_113_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_0_MPORT_113_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_0_MPORT_113_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_4_tile_v_3_MPORT_17_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_4_tile_v_3_MPORT_17_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_4_tile_v_3_MPORT_17_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_4_tile_v_2_MPORT_17_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_4_tile_v_2_MPORT_17_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_4_tile_v_2_MPORT_17_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_4_tile_v_1_MPORT_17_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_4_tile_v_1_MPORT_17_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_4_tile_v_1_MPORT_17_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_4_tile_v_0_MPORT_17_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_4_tile_v_0_MPORT_17_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_4_tile_v_0_MPORT_17_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_4_tile_v_3_MPORT_17_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_4_tile_v_3_MPORT_17_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_4_tile_v_3_MPORT_17_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_4_tile_v_2_MPORT_17_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_4_tile_v_2_MPORT_17_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_4_tile_v_2_MPORT_17_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_4_tile_v_1_MPORT_17_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_4_tile_v_1_MPORT_17_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_4_tile_v_1_MPORT_17_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_4_tile_v_0_MPORT_17_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_4_tile_v_0_MPORT_17_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_4_tile_v_0_MPORT_17_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_1_MPORT_114_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_1_MPORT_114_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_1_MPORT_114_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_0_MPORT_114_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_0_MPORT_114_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_0_MPORT_114_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_4_tile_v_3_MPORT_18_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_4_tile_v_3_MPORT_18_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_4_tile_v_3_MPORT_18_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_4_tile_v_2_MPORT_18_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_4_tile_v_2_MPORT_18_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_4_tile_v_2_MPORT_18_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_4_tile_v_1_MPORT_18_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_4_tile_v_1_MPORT_18_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_4_tile_v_1_MPORT_18_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_4_tile_v_0_MPORT_18_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_4_tile_v_0_MPORT_18_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_4_tile_v_0_MPORT_18_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_4_tile_v_3_MPORT_18_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_4_tile_v_3_MPORT_18_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_4_tile_v_3_MPORT_18_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_4_tile_v_2_MPORT_18_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_4_tile_v_2_MPORT_18_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_4_tile_v_2_MPORT_18_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_4_tile_v_1_MPORT_18_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_4_tile_v_1_MPORT_18_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_4_tile_v_1_MPORT_18_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_4_tile_v_0_MPORT_18_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_4_tile_v_0_MPORT_18_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_4_tile_v_0_MPORT_18_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_3_MPORT_38_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_3_MPORT_38_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_3_MPORT_38_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_2_MPORT_38_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_2_MPORT_38_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_2_MPORT_38_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_1_MPORT_115_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_1_MPORT_115_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_1_MPORT_115_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_0_MPORT_115_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_0_MPORT_115_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_0_MPORT_115_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_4_tile_v_3_MPORT_19_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_4_tile_v_3_MPORT_19_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_4_tile_v_3_MPORT_19_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_4_tile_v_2_MPORT_19_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_4_tile_v_2_MPORT_19_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_4_tile_v_2_MPORT_19_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_4_tile_v_1_MPORT_19_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_4_tile_v_1_MPORT_19_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_4_tile_v_1_MPORT_19_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_4_tile_v_0_MPORT_19_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_4_tile_v_0_MPORT_19_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_4_tile_v_0_MPORT_19_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_4_tile_v_3_MPORT_19_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_4_tile_v_3_MPORT_19_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_4_tile_v_3_MPORT_19_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_4_tile_v_2_MPORT_19_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_4_tile_v_2_MPORT_19_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_4_tile_v_2_MPORT_19_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_4_tile_v_1_MPORT_19_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_4_tile_v_1_MPORT_19_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_4_tile_v_1_MPORT_19_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_4_tile_v_0_MPORT_19_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_4_tile_v_0_MPORT_19_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_4_tile_v_0_MPORT_19_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_1_MPORT_116_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_1_MPORT_116_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_1_MPORT_116_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_0_MPORT_116_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_0_MPORT_116_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_0_MPORT_116_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_4_tile_v_3_MPORT_20_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_4_tile_v_3_MPORT_20_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_4_tile_v_3_MPORT_20_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_4_tile_v_2_MPORT_20_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_4_tile_v_2_MPORT_20_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_4_tile_v_2_MPORT_20_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_4_tile_v_1_MPORT_20_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_4_tile_v_1_MPORT_20_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_4_tile_v_1_MPORT_20_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_4_tile_v_0_MPORT_20_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_4_tile_v_0_MPORT_20_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_4_tile_v_0_MPORT_20_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_4_tile_v_3_MPORT_20_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_4_tile_v_3_MPORT_20_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_4_tile_v_3_MPORT_20_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_4_tile_v_2_MPORT_20_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_4_tile_v_2_MPORT_20_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_4_tile_v_2_MPORT_20_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_4_tile_v_1_MPORT_20_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_4_tile_v_1_MPORT_20_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_4_tile_v_1_MPORT_20_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_4_tile_v_0_MPORT_20_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_4_tile_v_0_MPORT_20_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_4_tile_v_0_MPORT_20_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_3_MPORT_39_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_3_MPORT_39_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_3_MPORT_39_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_2_MPORT_39_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_2_MPORT_39_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_2_MPORT_39_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_1_MPORT_117_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_1_MPORT_117_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_1_MPORT_117_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_0_MPORT_117_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_0_MPORT_117_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_0_MPORT_117_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_4_tile_v_3_MPORT_21_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_4_tile_v_3_MPORT_21_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_4_tile_v_3_MPORT_21_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_4_tile_v_2_MPORT_21_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_4_tile_v_2_MPORT_21_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_4_tile_v_2_MPORT_21_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_4_tile_v_1_MPORT_21_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_4_tile_v_1_MPORT_21_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_4_tile_v_1_MPORT_21_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_4_tile_v_0_MPORT_21_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_4_tile_v_0_MPORT_21_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_4_tile_v_0_MPORT_21_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_4_tile_v_3_MPORT_21_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_4_tile_v_3_MPORT_21_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_4_tile_v_3_MPORT_21_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_4_tile_v_2_MPORT_21_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_4_tile_v_2_MPORT_21_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_4_tile_v_2_MPORT_21_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_4_tile_v_1_MPORT_21_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_4_tile_v_1_MPORT_21_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_4_tile_v_1_MPORT_21_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_4_tile_v_0_MPORT_21_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_4_tile_v_0_MPORT_21_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_4_tile_v_0_MPORT_21_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_1_MPORT_118_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_1_MPORT_118_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_1_MPORT_118_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_0_MPORT_118_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_0_MPORT_118_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_0_MPORT_118_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_4_tile_v_3_MPORT_22_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_4_tile_v_3_MPORT_22_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_4_tile_v_3_MPORT_22_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_4_tile_v_2_MPORT_22_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_4_tile_v_2_MPORT_22_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_4_tile_v_2_MPORT_22_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_4_tile_v_1_MPORT_22_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_4_tile_v_1_MPORT_22_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_4_tile_v_1_MPORT_22_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_4_tile_v_0_MPORT_22_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_4_tile_v_0_MPORT_22_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_4_tile_v_0_MPORT_22_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_4_tile_v_3_MPORT_22_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_4_tile_v_3_MPORT_22_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_4_tile_v_3_MPORT_22_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_4_tile_v_2_MPORT_22_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_4_tile_v_2_MPORT_22_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_4_tile_v_2_MPORT_22_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_4_tile_v_1_MPORT_22_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_4_tile_v_1_MPORT_22_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_4_tile_v_1_MPORT_22_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_4_tile_v_0_MPORT_22_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_4_tile_v_0_MPORT_22_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_4_tile_v_0_MPORT_22_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_1_MPORT_119_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_1_MPORT_119_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_1_MPORT_119_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_0_MPORT_119_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_0_MPORT_119_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_0_MPORT_119_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_4_tile_v_3_MPORT_23_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_4_tile_v_3_MPORT_23_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_4_tile_v_3_MPORT_23_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_4_tile_v_2_MPORT_23_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_4_tile_v_2_MPORT_23_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_4_tile_v_2_MPORT_23_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_4_tile_v_1_MPORT_23_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_4_tile_v_1_MPORT_23_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_4_tile_v_1_MPORT_23_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_4_tile_v_0_MPORT_23_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_4_tile_v_0_MPORT_23_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_4_tile_v_0_MPORT_23_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_4_tile_v_3_MPORT_23_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_4_tile_v_3_MPORT_23_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_4_tile_v_3_MPORT_23_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_4_tile_v_2_MPORT_23_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_4_tile_v_2_MPORT_23_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_4_tile_v_2_MPORT_23_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_4_tile_v_1_MPORT_23_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_4_tile_v_1_MPORT_23_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_4_tile_v_1_MPORT_23_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_4_tile_v_0_MPORT_23_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_4_tile_v_0_MPORT_23_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_4_tile_v_0_MPORT_23_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_1_MPORT_120_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_1_MPORT_120_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_1_MPORT_120_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_0_MPORT_120_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_0_MPORT_120_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_0_MPORT_120_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_5_tile_v_3_MPORT_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_5_tile_v_3_MPORT_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_5_tile_v_3_MPORT_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_5_tile_v_2_MPORT_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_5_tile_v_2_MPORT_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_5_tile_v_2_MPORT_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_5_tile_v_1_MPORT_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_5_tile_v_1_MPORT_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_5_tile_v_1_MPORT_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_5_tile_v_0_MPORT_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_5_tile_v_0_MPORT_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_5_tile_v_0_MPORT_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_5_tile_v_3_MPORT_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_5_tile_v_3_MPORT_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_5_tile_v_3_MPORT_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_5_tile_v_2_MPORT_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_5_tile_v_2_MPORT_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_5_tile_v_2_MPORT_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_5_tile_v_1_MPORT_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_5_tile_v_1_MPORT_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_5_tile_v_1_MPORT_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_5_tile_v_0_MPORT_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_5_tile_v_0_MPORT_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_5_tile_v_0_MPORT_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_3_MPORT_40_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_3_MPORT_40_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_3_MPORT_40_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_2_MPORT_40_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_2_MPORT_40_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_2_MPORT_40_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_1_MPORT_121_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_1_MPORT_121_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_1_MPORT_121_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_0_MPORT_121_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_0_MPORT_121_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_0_MPORT_121_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_5_tile_v_3_MPORT_1_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_5_tile_v_3_MPORT_1_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_5_tile_v_3_MPORT_1_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_5_tile_v_2_MPORT_1_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_5_tile_v_2_MPORT_1_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_5_tile_v_2_MPORT_1_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_5_tile_v_1_MPORT_1_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_5_tile_v_1_MPORT_1_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_5_tile_v_1_MPORT_1_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_5_tile_v_0_MPORT_1_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_5_tile_v_0_MPORT_1_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_5_tile_v_0_MPORT_1_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_5_tile_v_3_MPORT_1_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_5_tile_v_3_MPORT_1_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_5_tile_v_3_MPORT_1_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_5_tile_v_2_MPORT_1_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_5_tile_v_2_MPORT_1_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_5_tile_v_2_MPORT_1_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_5_tile_v_1_MPORT_1_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_5_tile_v_1_MPORT_1_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_5_tile_v_1_MPORT_1_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_5_tile_v_0_MPORT_1_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_5_tile_v_0_MPORT_1_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_5_tile_v_0_MPORT_1_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_1_MPORT_122_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_1_MPORT_122_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_1_MPORT_122_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_0_MPORT_122_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_0_MPORT_122_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_0_MPORT_122_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_5_tile_v_3_MPORT_2_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_5_tile_v_3_MPORT_2_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_5_tile_v_3_MPORT_2_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_5_tile_v_2_MPORT_2_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_5_tile_v_2_MPORT_2_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_5_tile_v_2_MPORT_2_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_5_tile_v_1_MPORT_2_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_5_tile_v_1_MPORT_2_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_5_tile_v_1_MPORT_2_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_5_tile_v_0_MPORT_2_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_5_tile_v_0_MPORT_2_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_5_tile_v_0_MPORT_2_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_5_tile_v_3_MPORT_2_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_5_tile_v_3_MPORT_2_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_5_tile_v_3_MPORT_2_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_5_tile_v_2_MPORT_2_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_5_tile_v_2_MPORT_2_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_5_tile_v_2_MPORT_2_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_5_tile_v_1_MPORT_2_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_5_tile_v_1_MPORT_2_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_5_tile_v_1_MPORT_2_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_5_tile_v_0_MPORT_2_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_5_tile_v_0_MPORT_2_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_5_tile_v_0_MPORT_2_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_3_MPORT_41_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_3_MPORT_41_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_3_MPORT_41_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_2_MPORT_41_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_2_MPORT_41_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_2_MPORT_41_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_1_MPORT_123_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_1_MPORT_123_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_1_MPORT_123_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_0_MPORT_123_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_0_MPORT_123_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_0_MPORT_123_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_5_tile_v_3_MPORT_3_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_5_tile_v_3_MPORT_3_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_5_tile_v_3_MPORT_3_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_5_tile_v_2_MPORT_3_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_5_tile_v_2_MPORT_3_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_5_tile_v_2_MPORT_3_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_5_tile_v_1_MPORT_3_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_5_tile_v_1_MPORT_3_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_5_tile_v_1_MPORT_3_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_5_tile_v_0_MPORT_3_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_5_tile_v_0_MPORT_3_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_5_tile_v_0_MPORT_3_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_5_tile_v_3_MPORT_3_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_5_tile_v_3_MPORT_3_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_5_tile_v_3_MPORT_3_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_5_tile_v_2_MPORT_3_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_5_tile_v_2_MPORT_3_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_5_tile_v_2_MPORT_3_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_5_tile_v_1_MPORT_3_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_5_tile_v_1_MPORT_3_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_5_tile_v_1_MPORT_3_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_5_tile_v_0_MPORT_3_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_5_tile_v_0_MPORT_3_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_5_tile_v_0_MPORT_3_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_1_MPORT_124_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_1_MPORT_124_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_1_MPORT_124_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_0_MPORT_124_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_0_MPORT_124_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_0_MPORT_124_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_5_tile_v_3_MPORT_4_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_5_tile_v_3_MPORT_4_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_5_tile_v_3_MPORT_4_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_5_tile_v_2_MPORT_4_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_5_tile_v_2_MPORT_4_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_5_tile_v_2_MPORT_4_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_5_tile_v_1_MPORT_4_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_5_tile_v_1_MPORT_4_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_5_tile_v_1_MPORT_4_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_5_tile_v_0_MPORT_4_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_5_tile_v_0_MPORT_4_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_5_tile_v_0_MPORT_4_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_5_tile_v_3_MPORT_4_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_5_tile_v_3_MPORT_4_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_5_tile_v_3_MPORT_4_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_5_tile_v_2_MPORT_4_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_5_tile_v_2_MPORT_4_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_5_tile_v_2_MPORT_4_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_5_tile_v_1_MPORT_4_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_5_tile_v_1_MPORT_4_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_5_tile_v_1_MPORT_4_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_5_tile_v_0_MPORT_4_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_5_tile_v_0_MPORT_4_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_5_tile_v_0_MPORT_4_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_1_MPORT_125_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_1_MPORT_125_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_1_MPORT_125_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_0_MPORT_125_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_0_MPORT_125_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_0_MPORT_125_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_5_tile_v_3_MPORT_5_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_5_tile_v_3_MPORT_5_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_5_tile_v_3_MPORT_5_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_5_tile_v_2_MPORT_5_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_5_tile_v_2_MPORT_5_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_5_tile_v_2_MPORT_5_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_5_tile_v_1_MPORT_5_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_5_tile_v_1_MPORT_5_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_5_tile_v_1_MPORT_5_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_5_tile_v_0_MPORT_5_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_5_tile_v_0_MPORT_5_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_5_tile_v_0_MPORT_5_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_5_tile_v_3_MPORT_5_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_5_tile_v_3_MPORT_5_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_5_tile_v_3_MPORT_5_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_5_tile_v_2_MPORT_5_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_5_tile_v_2_MPORT_5_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_5_tile_v_2_MPORT_5_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_5_tile_v_1_MPORT_5_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_5_tile_v_1_MPORT_5_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_5_tile_v_1_MPORT_5_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_5_tile_v_0_MPORT_5_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_5_tile_v_0_MPORT_5_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_5_tile_v_0_MPORT_5_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_1_MPORT_126_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_1_MPORT_126_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_1_MPORT_126_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_0_MPORT_126_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_0_MPORT_126_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_0_MPORT_126_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_5_tile_v_3_MPORT_6_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_5_tile_v_3_MPORT_6_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_5_tile_v_3_MPORT_6_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_5_tile_v_2_MPORT_6_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_5_tile_v_2_MPORT_6_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_5_tile_v_2_MPORT_6_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_5_tile_v_1_MPORT_6_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_5_tile_v_1_MPORT_6_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_5_tile_v_1_MPORT_6_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_5_tile_v_0_MPORT_6_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_5_tile_v_0_MPORT_6_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_5_tile_v_0_MPORT_6_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_5_tile_v_3_MPORT_6_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_5_tile_v_3_MPORT_6_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_5_tile_v_3_MPORT_6_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_5_tile_v_2_MPORT_6_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_5_tile_v_2_MPORT_6_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_5_tile_v_2_MPORT_6_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_5_tile_v_1_MPORT_6_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_5_tile_v_1_MPORT_6_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_5_tile_v_1_MPORT_6_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_5_tile_v_0_MPORT_6_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_5_tile_v_0_MPORT_6_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_5_tile_v_0_MPORT_6_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_3_MPORT_42_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_3_MPORT_42_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_3_MPORT_42_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_2_MPORT_42_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_2_MPORT_42_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_2_MPORT_42_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_1_MPORT_127_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_1_MPORT_127_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_1_MPORT_127_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_0_MPORT_127_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_0_MPORT_127_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_0_MPORT_127_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_5_tile_v_3_MPORT_7_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_5_tile_v_3_MPORT_7_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_5_tile_v_3_MPORT_7_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_5_tile_v_2_MPORT_7_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_5_tile_v_2_MPORT_7_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_5_tile_v_2_MPORT_7_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_5_tile_v_1_MPORT_7_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_5_tile_v_1_MPORT_7_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_5_tile_v_1_MPORT_7_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_5_tile_v_0_MPORT_7_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_5_tile_v_0_MPORT_7_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_5_tile_v_0_MPORT_7_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_5_tile_v_3_MPORT_7_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_5_tile_v_3_MPORT_7_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_5_tile_v_3_MPORT_7_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_5_tile_v_2_MPORT_7_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_5_tile_v_2_MPORT_7_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_5_tile_v_2_MPORT_7_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_5_tile_v_1_MPORT_7_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_5_tile_v_1_MPORT_7_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_5_tile_v_1_MPORT_7_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_5_tile_v_0_MPORT_7_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_5_tile_v_0_MPORT_7_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_5_tile_v_0_MPORT_7_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_1_MPORT_128_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_1_MPORT_128_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_1_MPORT_128_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_0_MPORT_128_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_0_MPORT_128_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_0_MPORT_128_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_5_tile_v_3_MPORT_8_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_5_tile_v_3_MPORT_8_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_5_tile_v_3_MPORT_8_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_5_tile_v_2_MPORT_8_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_5_tile_v_2_MPORT_8_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_5_tile_v_2_MPORT_8_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_5_tile_v_1_MPORT_8_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_5_tile_v_1_MPORT_8_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_5_tile_v_1_MPORT_8_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_5_tile_v_0_MPORT_8_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_5_tile_v_0_MPORT_8_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_5_tile_v_0_MPORT_8_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_5_tile_v_3_MPORT_8_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_5_tile_v_3_MPORT_8_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_5_tile_v_3_MPORT_8_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_5_tile_v_2_MPORT_8_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_5_tile_v_2_MPORT_8_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_5_tile_v_2_MPORT_8_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_5_tile_v_1_MPORT_8_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_5_tile_v_1_MPORT_8_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_5_tile_v_1_MPORT_8_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_5_tile_v_0_MPORT_8_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_5_tile_v_0_MPORT_8_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_5_tile_v_0_MPORT_8_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_3_MPORT_43_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_3_MPORT_43_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_3_MPORT_43_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_2_MPORT_43_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_2_MPORT_43_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_2_MPORT_43_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_1_MPORT_129_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_1_MPORT_129_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_1_MPORT_129_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_0_MPORT_129_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_0_MPORT_129_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_0_MPORT_129_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_5_tile_v_3_MPORT_9_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_5_tile_v_3_MPORT_9_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_5_tile_v_3_MPORT_9_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_5_tile_v_2_MPORT_9_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_5_tile_v_2_MPORT_9_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_5_tile_v_2_MPORT_9_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_5_tile_v_1_MPORT_9_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_5_tile_v_1_MPORT_9_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_5_tile_v_1_MPORT_9_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_5_tile_v_0_MPORT_9_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_5_tile_v_0_MPORT_9_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_5_tile_v_0_MPORT_9_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_5_tile_v_3_MPORT_9_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_5_tile_v_3_MPORT_9_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_5_tile_v_3_MPORT_9_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_5_tile_v_2_MPORT_9_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_5_tile_v_2_MPORT_9_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_5_tile_v_2_MPORT_9_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_5_tile_v_1_MPORT_9_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_5_tile_v_1_MPORT_9_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_5_tile_v_1_MPORT_9_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_5_tile_v_0_MPORT_9_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_5_tile_v_0_MPORT_9_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_5_tile_v_0_MPORT_9_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_1_MPORT_130_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_1_MPORT_130_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_1_MPORT_130_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_0_MPORT_130_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_0_MPORT_130_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_0_MPORT_130_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_5_tile_v_3_MPORT_10_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_5_tile_v_3_MPORT_10_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_5_tile_v_3_MPORT_10_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_5_tile_v_2_MPORT_10_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_5_tile_v_2_MPORT_10_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_5_tile_v_2_MPORT_10_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_5_tile_v_1_MPORT_10_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_5_tile_v_1_MPORT_10_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_5_tile_v_1_MPORT_10_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_5_tile_v_0_MPORT_10_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_5_tile_v_0_MPORT_10_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_5_tile_v_0_MPORT_10_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_5_tile_v_3_MPORT_10_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_5_tile_v_3_MPORT_10_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_5_tile_v_3_MPORT_10_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_5_tile_v_2_MPORT_10_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_5_tile_v_2_MPORT_10_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_5_tile_v_2_MPORT_10_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_5_tile_v_1_MPORT_10_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_5_tile_v_1_MPORT_10_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_5_tile_v_1_MPORT_10_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_5_tile_v_0_MPORT_10_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_5_tile_v_0_MPORT_10_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_5_tile_v_0_MPORT_10_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_1_MPORT_131_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_1_MPORT_131_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_1_MPORT_131_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_0_MPORT_131_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_0_MPORT_131_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_0_MPORT_131_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_5_tile_v_3_MPORT_11_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_5_tile_v_3_MPORT_11_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_5_tile_v_3_MPORT_11_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_5_tile_v_2_MPORT_11_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_5_tile_v_2_MPORT_11_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_5_tile_v_2_MPORT_11_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_5_tile_v_1_MPORT_11_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_5_tile_v_1_MPORT_11_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_5_tile_v_1_MPORT_11_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_5_tile_v_0_MPORT_11_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_5_tile_v_0_MPORT_11_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_5_tile_v_0_MPORT_11_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_5_tile_v_3_MPORT_11_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_5_tile_v_3_MPORT_11_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_5_tile_v_3_MPORT_11_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_5_tile_v_2_MPORT_11_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_5_tile_v_2_MPORT_11_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_5_tile_v_2_MPORT_11_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_5_tile_v_1_MPORT_11_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_5_tile_v_1_MPORT_11_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_5_tile_v_1_MPORT_11_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_5_tile_v_0_MPORT_11_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_5_tile_v_0_MPORT_11_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_5_tile_v_0_MPORT_11_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_1_MPORT_132_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_1_MPORT_132_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_1_MPORT_132_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_0_MPORT_132_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_0_MPORT_132_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_0_MPORT_132_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_5_tile_v_3_MPORT_12_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_5_tile_v_3_MPORT_12_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_5_tile_v_3_MPORT_12_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_5_tile_v_2_MPORT_12_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_5_tile_v_2_MPORT_12_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_5_tile_v_2_MPORT_12_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_5_tile_v_1_MPORT_12_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_5_tile_v_1_MPORT_12_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_5_tile_v_1_MPORT_12_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_5_tile_v_0_MPORT_12_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_5_tile_v_0_MPORT_12_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_5_tile_v_0_MPORT_12_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_5_tile_v_3_MPORT_12_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_5_tile_v_3_MPORT_12_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_5_tile_v_3_MPORT_12_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_5_tile_v_2_MPORT_12_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_5_tile_v_2_MPORT_12_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_5_tile_v_2_MPORT_12_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_5_tile_v_1_MPORT_12_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_5_tile_v_1_MPORT_12_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_5_tile_v_1_MPORT_12_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_5_tile_v_0_MPORT_12_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_5_tile_v_0_MPORT_12_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_5_tile_v_0_MPORT_12_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_3_MPORT_44_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_3_MPORT_44_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_3_MPORT_44_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_2_MPORT_44_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_2_MPORT_44_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_2_MPORT_44_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_1_MPORT_133_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_1_MPORT_133_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_1_MPORT_133_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_0_MPORT_133_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_0_MPORT_133_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_0_MPORT_133_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_5_tile_v_3_MPORT_13_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_5_tile_v_3_MPORT_13_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_5_tile_v_3_MPORT_13_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_5_tile_v_2_MPORT_13_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_5_tile_v_2_MPORT_13_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_5_tile_v_2_MPORT_13_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_5_tile_v_1_MPORT_13_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_5_tile_v_1_MPORT_13_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_5_tile_v_1_MPORT_13_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_5_tile_v_0_MPORT_13_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_5_tile_v_0_MPORT_13_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_5_tile_v_0_MPORT_13_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_5_tile_v_3_MPORT_13_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_5_tile_v_3_MPORT_13_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_5_tile_v_3_MPORT_13_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_5_tile_v_2_MPORT_13_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_5_tile_v_2_MPORT_13_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_5_tile_v_2_MPORT_13_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_5_tile_v_1_MPORT_13_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_5_tile_v_1_MPORT_13_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_5_tile_v_1_MPORT_13_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_5_tile_v_0_MPORT_13_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_5_tile_v_0_MPORT_13_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_5_tile_v_0_MPORT_13_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_1_MPORT_134_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_1_MPORT_134_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_1_MPORT_134_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_0_MPORT_134_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_0_MPORT_134_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_0_MPORT_134_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_5_tile_v_3_MPORT_14_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_5_tile_v_3_MPORT_14_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_5_tile_v_3_MPORT_14_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_5_tile_v_2_MPORT_14_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_5_tile_v_2_MPORT_14_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_5_tile_v_2_MPORT_14_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_5_tile_v_1_MPORT_14_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_5_tile_v_1_MPORT_14_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_5_tile_v_1_MPORT_14_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_5_tile_v_0_MPORT_14_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_5_tile_v_0_MPORT_14_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_5_tile_v_0_MPORT_14_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_5_tile_v_3_MPORT_14_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_5_tile_v_3_MPORT_14_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_5_tile_v_3_MPORT_14_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_5_tile_v_2_MPORT_14_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_5_tile_v_2_MPORT_14_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_5_tile_v_2_MPORT_14_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_5_tile_v_1_MPORT_14_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_5_tile_v_1_MPORT_14_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_5_tile_v_1_MPORT_14_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_5_tile_v_0_MPORT_14_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_5_tile_v_0_MPORT_14_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_5_tile_v_0_MPORT_14_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_3_MPORT_45_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_3_MPORT_45_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_3_MPORT_45_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_2_MPORT_45_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_2_MPORT_45_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_2_MPORT_45_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_1_MPORT_135_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_1_MPORT_135_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_1_MPORT_135_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_0_MPORT_135_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_0_MPORT_135_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_0_MPORT_135_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_5_tile_v_3_MPORT_15_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_5_tile_v_3_MPORT_15_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_5_tile_v_3_MPORT_15_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_5_tile_v_2_MPORT_15_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_5_tile_v_2_MPORT_15_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_5_tile_v_2_MPORT_15_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_5_tile_v_1_MPORT_15_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_5_tile_v_1_MPORT_15_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_5_tile_v_1_MPORT_15_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_5_tile_v_0_MPORT_15_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_5_tile_v_0_MPORT_15_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_5_tile_v_0_MPORT_15_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_5_tile_v_3_MPORT_15_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_5_tile_v_3_MPORT_15_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_5_tile_v_3_MPORT_15_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_5_tile_v_2_MPORT_15_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_5_tile_v_2_MPORT_15_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_5_tile_v_2_MPORT_15_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_5_tile_v_1_MPORT_15_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_5_tile_v_1_MPORT_15_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_5_tile_v_1_MPORT_15_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_5_tile_v_0_MPORT_15_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_5_tile_v_0_MPORT_15_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_5_tile_v_0_MPORT_15_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_1_MPORT_136_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_1_MPORT_136_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_1_MPORT_136_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_0_MPORT_136_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_0_MPORT_136_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_0_MPORT_136_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_5_tile_v_3_MPORT_16_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_5_tile_v_3_MPORT_16_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_5_tile_v_3_MPORT_16_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_5_tile_v_2_MPORT_16_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_5_tile_v_2_MPORT_16_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_5_tile_v_2_MPORT_16_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_5_tile_v_1_MPORT_16_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_5_tile_v_1_MPORT_16_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_5_tile_v_1_MPORT_16_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_5_tile_v_0_MPORT_16_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_5_tile_v_0_MPORT_16_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_5_tile_v_0_MPORT_16_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_5_tile_v_3_MPORT_16_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_5_tile_v_3_MPORT_16_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_5_tile_v_3_MPORT_16_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_5_tile_v_2_MPORT_16_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_5_tile_v_2_MPORT_16_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_5_tile_v_2_MPORT_16_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_5_tile_v_1_MPORT_16_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_5_tile_v_1_MPORT_16_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_5_tile_v_1_MPORT_16_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_5_tile_v_0_MPORT_16_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_5_tile_v_0_MPORT_16_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_5_tile_v_0_MPORT_16_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_1_MPORT_137_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_1_MPORT_137_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_1_MPORT_137_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_0_MPORT_137_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_0_MPORT_137_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_0_MPORT_137_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_5_tile_v_3_MPORT_17_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_5_tile_v_3_MPORT_17_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_5_tile_v_3_MPORT_17_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_5_tile_v_2_MPORT_17_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_5_tile_v_2_MPORT_17_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_5_tile_v_2_MPORT_17_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_5_tile_v_1_MPORT_17_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_5_tile_v_1_MPORT_17_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_5_tile_v_1_MPORT_17_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_5_tile_v_0_MPORT_17_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_5_tile_v_0_MPORT_17_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_5_tile_v_0_MPORT_17_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_5_tile_v_3_MPORT_17_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_5_tile_v_3_MPORT_17_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_5_tile_v_3_MPORT_17_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_5_tile_v_2_MPORT_17_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_5_tile_v_2_MPORT_17_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_5_tile_v_2_MPORT_17_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_5_tile_v_1_MPORT_17_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_5_tile_v_1_MPORT_17_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_5_tile_v_1_MPORT_17_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_5_tile_v_0_MPORT_17_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_5_tile_v_0_MPORT_17_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_5_tile_v_0_MPORT_17_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_1_MPORT_138_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_1_MPORT_138_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_1_MPORT_138_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_0_MPORT_138_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_0_MPORT_138_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_0_MPORT_138_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_5_tile_v_3_MPORT_18_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_5_tile_v_3_MPORT_18_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_5_tile_v_3_MPORT_18_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_5_tile_v_2_MPORT_18_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_5_tile_v_2_MPORT_18_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_5_tile_v_2_MPORT_18_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_5_tile_v_1_MPORT_18_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_5_tile_v_1_MPORT_18_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_5_tile_v_1_MPORT_18_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_5_tile_v_0_MPORT_18_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_5_tile_v_0_MPORT_18_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_5_tile_v_0_MPORT_18_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_5_tile_v_3_MPORT_18_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_5_tile_v_3_MPORT_18_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_5_tile_v_3_MPORT_18_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_5_tile_v_2_MPORT_18_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_5_tile_v_2_MPORT_18_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_5_tile_v_2_MPORT_18_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_5_tile_v_1_MPORT_18_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_5_tile_v_1_MPORT_18_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_5_tile_v_1_MPORT_18_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_5_tile_v_0_MPORT_18_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_5_tile_v_0_MPORT_18_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_5_tile_v_0_MPORT_18_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_3_MPORT_46_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_3_MPORT_46_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_3_MPORT_46_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_2_MPORT_46_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_2_MPORT_46_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_2_MPORT_46_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_1_MPORT_139_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_1_MPORT_139_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_1_MPORT_139_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_0_MPORT_139_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_0_MPORT_139_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_0_MPORT_139_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_5_tile_v_3_MPORT_19_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_5_tile_v_3_MPORT_19_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_5_tile_v_3_MPORT_19_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_5_tile_v_2_MPORT_19_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_5_tile_v_2_MPORT_19_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_5_tile_v_2_MPORT_19_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_5_tile_v_1_MPORT_19_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_5_tile_v_1_MPORT_19_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_5_tile_v_1_MPORT_19_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_5_tile_v_0_MPORT_19_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_5_tile_v_0_MPORT_19_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_5_tile_v_0_MPORT_19_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_5_tile_v_3_MPORT_19_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_5_tile_v_3_MPORT_19_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_5_tile_v_3_MPORT_19_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_5_tile_v_2_MPORT_19_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_5_tile_v_2_MPORT_19_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_5_tile_v_2_MPORT_19_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_5_tile_v_1_MPORT_19_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_5_tile_v_1_MPORT_19_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_5_tile_v_1_MPORT_19_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_5_tile_v_0_MPORT_19_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_5_tile_v_0_MPORT_19_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_5_tile_v_0_MPORT_19_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_1_MPORT_140_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_1_MPORT_140_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_1_MPORT_140_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_0_MPORT_140_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_0_MPORT_140_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_0_MPORT_140_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_5_tile_v_3_MPORT_20_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_5_tile_v_3_MPORT_20_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_5_tile_v_3_MPORT_20_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_5_tile_v_2_MPORT_20_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_5_tile_v_2_MPORT_20_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_5_tile_v_2_MPORT_20_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_5_tile_v_1_MPORT_20_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_5_tile_v_1_MPORT_20_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_5_tile_v_1_MPORT_20_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_5_tile_v_0_MPORT_20_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_5_tile_v_0_MPORT_20_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_5_tile_v_0_MPORT_20_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_5_tile_v_3_MPORT_20_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_5_tile_v_3_MPORT_20_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_5_tile_v_3_MPORT_20_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_5_tile_v_2_MPORT_20_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_5_tile_v_2_MPORT_20_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_5_tile_v_2_MPORT_20_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_5_tile_v_1_MPORT_20_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_5_tile_v_1_MPORT_20_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_5_tile_v_1_MPORT_20_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_5_tile_v_0_MPORT_20_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_5_tile_v_0_MPORT_20_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_5_tile_v_0_MPORT_20_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_3_MPORT_47_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_3_MPORT_47_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_3_MPORT_47_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_2_MPORT_47_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_2_MPORT_47_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_2_MPORT_47_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_1_MPORT_141_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_1_MPORT_141_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_1_MPORT_141_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_0_MPORT_141_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_0_MPORT_141_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_0_MPORT_141_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_5_tile_v_3_MPORT_21_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_5_tile_v_3_MPORT_21_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_5_tile_v_3_MPORT_21_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_5_tile_v_2_MPORT_21_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_5_tile_v_2_MPORT_21_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_5_tile_v_2_MPORT_21_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_5_tile_v_1_MPORT_21_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_5_tile_v_1_MPORT_21_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_5_tile_v_1_MPORT_21_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_5_tile_v_0_MPORT_21_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_5_tile_v_0_MPORT_21_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_5_tile_v_0_MPORT_21_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_5_tile_v_3_MPORT_21_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_5_tile_v_3_MPORT_21_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_5_tile_v_3_MPORT_21_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_5_tile_v_2_MPORT_21_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_5_tile_v_2_MPORT_21_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_5_tile_v_2_MPORT_21_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_5_tile_v_1_MPORT_21_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_5_tile_v_1_MPORT_21_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_5_tile_v_1_MPORT_21_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_5_tile_v_0_MPORT_21_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_5_tile_v_0_MPORT_21_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_5_tile_v_0_MPORT_21_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_1_MPORT_142_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_1_MPORT_142_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_1_MPORT_142_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_0_MPORT_142_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_0_MPORT_142_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_0_MPORT_142_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_5_tile_v_3_MPORT_22_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_5_tile_v_3_MPORT_22_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_5_tile_v_3_MPORT_22_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_5_tile_v_2_MPORT_22_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_5_tile_v_2_MPORT_22_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_5_tile_v_2_MPORT_22_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_5_tile_v_1_MPORT_22_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_5_tile_v_1_MPORT_22_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_5_tile_v_1_MPORT_22_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_5_tile_v_0_MPORT_22_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_5_tile_v_0_MPORT_22_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_5_tile_v_0_MPORT_22_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_5_tile_v_3_MPORT_22_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_5_tile_v_3_MPORT_22_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_5_tile_v_3_MPORT_22_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_5_tile_v_2_MPORT_22_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_5_tile_v_2_MPORT_22_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_5_tile_v_2_MPORT_22_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_5_tile_v_1_MPORT_22_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_5_tile_v_1_MPORT_22_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_5_tile_v_1_MPORT_22_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_5_tile_v_0_MPORT_22_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_5_tile_v_0_MPORT_22_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_5_tile_v_0_MPORT_22_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_1_MPORT_143_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_1_MPORT_143_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_1_MPORT_143_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_0_MPORT_143_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_0_MPORT_143_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_0_MPORT_143_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_5_tile_v_3_MPORT_23_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_5_tile_v_3_MPORT_23_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_5_tile_v_3_MPORT_23_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_5_tile_v_2_MPORT_23_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_5_tile_v_2_MPORT_23_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_5_tile_v_2_MPORT_23_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_5_tile_v_1_MPORT_23_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_5_tile_v_1_MPORT_23_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_5_tile_v_1_MPORT_23_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_5_tile_v_0_MPORT_23_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_5_tile_v_0_MPORT_23_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_5_tile_v_0_MPORT_23_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_5_tile_v_3_MPORT_23_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_5_tile_v_3_MPORT_23_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_5_tile_v_3_MPORT_23_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_5_tile_v_2_MPORT_23_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_5_tile_v_2_MPORT_23_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_5_tile_v_2_MPORT_23_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_5_tile_v_1_MPORT_23_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_5_tile_v_1_MPORT_23_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_5_tile_v_1_MPORT_23_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_5_tile_v_0_MPORT_23_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_5_tile_v_0_MPORT_23_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_5_tile_v_0_MPORT_23_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_1_MPORT_144_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_1_MPORT_144_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_1_MPORT_144_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_0_MPORT_144_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_0_MPORT_144_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_0_MPORT_144_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_6_tile_v_3_MPORT_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_6_tile_v_3_MPORT_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_6_tile_v_3_MPORT_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_6_tile_v_2_MPORT_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_6_tile_v_2_MPORT_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_6_tile_v_2_MPORT_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_6_tile_v_1_MPORT_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_6_tile_v_1_MPORT_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_6_tile_v_1_MPORT_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_6_tile_v_0_MPORT_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_6_tile_v_0_MPORT_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_6_tile_v_0_MPORT_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_6_tile_v_3_MPORT_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_6_tile_v_3_MPORT_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_6_tile_v_3_MPORT_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_6_tile_v_2_MPORT_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_6_tile_v_2_MPORT_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_6_tile_v_2_MPORT_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_6_tile_v_1_MPORT_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_6_tile_v_1_MPORT_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_6_tile_v_1_MPORT_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_6_tile_v_0_MPORT_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_6_tile_v_0_MPORT_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_6_tile_v_0_MPORT_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_3_MPORT_48_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_3_MPORT_48_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_3_MPORT_48_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_2_MPORT_48_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_2_MPORT_48_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_2_MPORT_48_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_1_MPORT_145_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_1_MPORT_145_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_1_MPORT_145_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_0_MPORT_145_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_0_MPORT_145_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_0_MPORT_145_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_6_tile_v_3_MPORT_1_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_6_tile_v_3_MPORT_1_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_6_tile_v_3_MPORT_1_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_6_tile_v_2_MPORT_1_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_6_tile_v_2_MPORT_1_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_6_tile_v_2_MPORT_1_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_6_tile_v_1_MPORT_1_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_6_tile_v_1_MPORT_1_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_6_tile_v_1_MPORT_1_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_6_tile_v_0_MPORT_1_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_6_tile_v_0_MPORT_1_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_6_tile_v_0_MPORT_1_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_6_tile_v_3_MPORT_1_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_6_tile_v_3_MPORT_1_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_6_tile_v_3_MPORT_1_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_6_tile_v_2_MPORT_1_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_6_tile_v_2_MPORT_1_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_6_tile_v_2_MPORT_1_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_6_tile_v_1_MPORT_1_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_6_tile_v_1_MPORT_1_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_6_tile_v_1_MPORT_1_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_6_tile_v_0_MPORT_1_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_6_tile_v_0_MPORT_1_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_6_tile_v_0_MPORT_1_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_1_MPORT_146_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_1_MPORT_146_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_1_MPORT_146_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_0_MPORT_146_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_0_MPORT_146_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_0_MPORT_146_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_6_tile_v_3_MPORT_2_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_6_tile_v_3_MPORT_2_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_6_tile_v_3_MPORT_2_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_6_tile_v_2_MPORT_2_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_6_tile_v_2_MPORT_2_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_6_tile_v_2_MPORT_2_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_6_tile_v_1_MPORT_2_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_6_tile_v_1_MPORT_2_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_6_tile_v_1_MPORT_2_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_6_tile_v_0_MPORT_2_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_6_tile_v_0_MPORT_2_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_6_tile_v_0_MPORT_2_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_6_tile_v_3_MPORT_2_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_6_tile_v_3_MPORT_2_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_6_tile_v_3_MPORT_2_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_6_tile_v_2_MPORT_2_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_6_tile_v_2_MPORT_2_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_6_tile_v_2_MPORT_2_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_6_tile_v_1_MPORT_2_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_6_tile_v_1_MPORT_2_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_6_tile_v_1_MPORT_2_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_6_tile_v_0_MPORT_2_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_6_tile_v_0_MPORT_2_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_6_tile_v_0_MPORT_2_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_3_MPORT_49_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_3_MPORT_49_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_3_MPORT_49_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_2_MPORT_49_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_2_MPORT_49_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_2_MPORT_49_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_1_MPORT_147_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_1_MPORT_147_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_1_MPORT_147_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_0_MPORT_147_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_0_MPORT_147_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_0_MPORT_147_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_6_tile_v_3_MPORT_3_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_6_tile_v_3_MPORT_3_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_6_tile_v_3_MPORT_3_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_6_tile_v_2_MPORT_3_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_6_tile_v_2_MPORT_3_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_6_tile_v_2_MPORT_3_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_6_tile_v_1_MPORT_3_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_6_tile_v_1_MPORT_3_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_6_tile_v_1_MPORT_3_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_6_tile_v_0_MPORT_3_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_6_tile_v_0_MPORT_3_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_6_tile_v_0_MPORT_3_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_6_tile_v_3_MPORT_3_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_6_tile_v_3_MPORT_3_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_6_tile_v_3_MPORT_3_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_6_tile_v_2_MPORT_3_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_6_tile_v_2_MPORT_3_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_6_tile_v_2_MPORT_3_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_6_tile_v_1_MPORT_3_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_6_tile_v_1_MPORT_3_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_6_tile_v_1_MPORT_3_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_6_tile_v_0_MPORT_3_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_6_tile_v_0_MPORT_3_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_6_tile_v_0_MPORT_3_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_1_MPORT_148_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_1_MPORT_148_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_1_MPORT_148_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_0_MPORT_148_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_0_MPORT_148_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_0_MPORT_148_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_6_tile_v_3_MPORT_4_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_6_tile_v_3_MPORT_4_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_6_tile_v_3_MPORT_4_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_6_tile_v_2_MPORT_4_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_6_tile_v_2_MPORT_4_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_6_tile_v_2_MPORT_4_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_6_tile_v_1_MPORT_4_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_6_tile_v_1_MPORT_4_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_6_tile_v_1_MPORT_4_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_6_tile_v_0_MPORT_4_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_6_tile_v_0_MPORT_4_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_6_tile_v_0_MPORT_4_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_6_tile_v_3_MPORT_4_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_6_tile_v_3_MPORT_4_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_6_tile_v_3_MPORT_4_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_6_tile_v_2_MPORT_4_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_6_tile_v_2_MPORT_4_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_6_tile_v_2_MPORT_4_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_6_tile_v_1_MPORT_4_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_6_tile_v_1_MPORT_4_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_6_tile_v_1_MPORT_4_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_6_tile_v_0_MPORT_4_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_6_tile_v_0_MPORT_4_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_6_tile_v_0_MPORT_4_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_1_MPORT_149_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_1_MPORT_149_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_1_MPORT_149_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_0_MPORT_149_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_0_MPORT_149_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_0_MPORT_149_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_6_tile_v_3_MPORT_5_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_6_tile_v_3_MPORT_5_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_6_tile_v_3_MPORT_5_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_6_tile_v_2_MPORT_5_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_6_tile_v_2_MPORT_5_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_6_tile_v_2_MPORT_5_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_6_tile_v_1_MPORT_5_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_6_tile_v_1_MPORT_5_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_6_tile_v_1_MPORT_5_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_6_tile_v_0_MPORT_5_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_6_tile_v_0_MPORT_5_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_6_tile_v_0_MPORT_5_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_6_tile_v_3_MPORT_5_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_6_tile_v_3_MPORT_5_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_6_tile_v_3_MPORT_5_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_6_tile_v_2_MPORT_5_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_6_tile_v_2_MPORT_5_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_6_tile_v_2_MPORT_5_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_6_tile_v_1_MPORT_5_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_6_tile_v_1_MPORT_5_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_6_tile_v_1_MPORT_5_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_6_tile_v_0_MPORT_5_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_6_tile_v_0_MPORT_5_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_6_tile_v_0_MPORT_5_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_1_MPORT_150_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_1_MPORT_150_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_1_MPORT_150_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_0_MPORT_150_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_0_MPORT_150_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_0_MPORT_150_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_6_tile_v_3_MPORT_6_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_6_tile_v_3_MPORT_6_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_6_tile_v_3_MPORT_6_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_6_tile_v_2_MPORT_6_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_6_tile_v_2_MPORT_6_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_6_tile_v_2_MPORT_6_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_6_tile_v_1_MPORT_6_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_6_tile_v_1_MPORT_6_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_6_tile_v_1_MPORT_6_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_6_tile_v_0_MPORT_6_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_6_tile_v_0_MPORT_6_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_6_tile_v_0_MPORT_6_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_6_tile_v_3_MPORT_6_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_6_tile_v_3_MPORT_6_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_6_tile_v_3_MPORT_6_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_6_tile_v_2_MPORT_6_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_6_tile_v_2_MPORT_6_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_6_tile_v_2_MPORT_6_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_6_tile_v_1_MPORT_6_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_6_tile_v_1_MPORT_6_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_6_tile_v_1_MPORT_6_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_6_tile_v_0_MPORT_6_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_6_tile_v_0_MPORT_6_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_6_tile_v_0_MPORT_6_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_3_MPORT_50_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_3_MPORT_50_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_3_MPORT_50_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_2_MPORT_50_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_2_MPORT_50_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_2_MPORT_50_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_1_MPORT_151_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_1_MPORT_151_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_1_MPORT_151_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_0_MPORT_151_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_0_MPORT_151_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_0_MPORT_151_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_6_tile_v_3_MPORT_7_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_6_tile_v_3_MPORT_7_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_6_tile_v_3_MPORT_7_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_6_tile_v_2_MPORT_7_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_6_tile_v_2_MPORT_7_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_6_tile_v_2_MPORT_7_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_6_tile_v_1_MPORT_7_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_6_tile_v_1_MPORT_7_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_6_tile_v_1_MPORT_7_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_6_tile_v_0_MPORT_7_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_6_tile_v_0_MPORT_7_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_6_tile_v_0_MPORT_7_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_6_tile_v_3_MPORT_7_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_6_tile_v_3_MPORT_7_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_6_tile_v_3_MPORT_7_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_6_tile_v_2_MPORT_7_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_6_tile_v_2_MPORT_7_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_6_tile_v_2_MPORT_7_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_6_tile_v_1_MPORT_7_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_6_tile_v_1_MPORT_7_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_6_tile_v_1_MPORT_7_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_6_tile_v_0_MPORT_7_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_6_tile_v_0_MPORT_7_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_6_tile_v_0_MPORT_7_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_1_MPORT_152_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_1_MPORT_152_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_1_MPORT_152_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_0_MPORT_152_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_0_MPORT_152_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_0_MPORT_152_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_6_tile_v_3_MPORT_8_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_6_tile_v_3_MPORT_8_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_6_tile_v_3_MPORT_8_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_6_tile_v_2_MPORT_8_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_6_tile_v_2_MPORT_8_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_6_tile_v_2_MPORT_8_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_6_tile_v_1_MPORT_8_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_6_tile_v_1_MPORT_8_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_6_tile_v_1_MPORT_8_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_6_tile_v_0_MPORT_8_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_6_tile_v_0_MPORT_8_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_6_tile_v_0_MPORT_8_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_6_tile_v_3_MPORT_8_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_6_tile_v_3_MPORT_8_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_6_tile_v_3_MPORT_8_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_6_tile_v_2_MPORT_8_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_6_tile_v_2_MPORT_8_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_6_tile_v_2_MPORT_8_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_6_tile_v_1_MPORT_8_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_6_tile_v_1_MPORT_8_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_6_tile_v_1_MPORT_8_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_6_tile_v_0_MPORT_8_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_6_tile_v_0_MPORT_8_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_6_tile_v_0_MPORT_8_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_3_MPORT_51_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_3_MPORT_51_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_3_MPORT_51_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_2_MPORT_51_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_2_MPORT_51_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_2_MPORT_51_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_1_MPORT_153_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_1_MPORT_153_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_1_MPORT_153_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_0_MPORT_153_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_0_MPORT_153_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_0_MPORT_153_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_6_tile_v_3_MPORT_9_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_6_tile_v_3_MPORT_9_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_6_tile_v_3_MPORT_9_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_6_tile_v_2_MPORT_9_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_6_tile_v_2_MPORT_9_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_6_tile_v_2_MPORT_9_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_6_tile_v_1_MPORT_9_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_6_tile_v_1_MPORT_9_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_6_tile_v_1_MPORT_9_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_6_tile_v_0_MPORT_9_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_6_tile_v_0_MPORT_9_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_6_tile_v_0_MPORT_9_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_6_tile_v_3_MPORT_9_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_6_tile_v_3_MPORT_9_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_6_tile_v_3_MPORT_9_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_6_tile_v_2_MPORT_9_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_6_tile_v_2_MPORT_9_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_6_tile_v_2_MPORT_9_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_6_tile_v_1_MPORT_9_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_6_tile_v_1_MPORT_9_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_6_tile_v_1_MPORT_9_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_6_tile_v_0_MPORT_9_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_6_tile_v_0_MPORT_9_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_6_tile_v_0_MPORT_9_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_1_MPORT_154_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_1_MPORT_154_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_1_MPORT_154_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_0_MPORT_154_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_0_MPORT_154_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_0_MPORT_154_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_6_tile_v_3_MPORT_10_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_6_tile_v_3_MPORT_10_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_6_tile_v_3_MPORT_10_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_6_tile_v_2_MPORT_10_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_6_tile_v_2_MPORT_10_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_6_tile_v_2_MPORT_10_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_6_tile_v_1_MPORT_10_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_6_tile_v_1_MPORT_10_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_6_tile_v_1_MPORT_10_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_6_tile_v_0_MPORT_10_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_6_tile_v_0_MPORT_10_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_6_tile_v_0_MPORT_10_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_6_tile_v_3_MPORT_10_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_6_tile_v_3_MPORT_10_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_6_tile_v_3_MPORT_10_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_6_tile_v_2_MPORT_10_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_6_tile_v_2_MPORT_10_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_6_tile_v_2_MPORT_10_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_6_tile_v_1_MPORT_10_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_6_tile_v_1_MPORT_10_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_6_tile_v_1_MPORT_10_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_6_tile_v_0_MPORT_10_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_6_tile_v_0_MPORT_10_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_6_tile_v_0_MPORT_10_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_1_MPORT_155_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_1_MPORT_155_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_1_MPORT_155_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_0_MPORT_155_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_0_MPORT_155_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_0_MPORT_155_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_6_tile_v_3_MPORT_11_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_6_tile_v_3_MPORT_11_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_6_tile_v_3_MPORT_11_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_6_tile_v_2_MPORT_11_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_6_tile_v_2_MPORT_11_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_6_tile_v_2_MPORT_11_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_6_tile_v_1_MPORT_11_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_6_tile_v_1_MPORT_11_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_6_tile_v_1_MPORT_11_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_6_tile_v_0_MPORT_11_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_6_tile_v_0_MPORT_11_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_6_tile_v_0_MPORT_11_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_6_tile_v_3_MPORT_11_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_6_tile_v_3_MPORT_11_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_6_tile_v_3_MPORT_11_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_6_tile_v_2_MPORT_11_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_6_tile_v_2_MPORT_11_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_6_tile_v_2_MPORT_11_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_6_tile_v_1_MPORT_11_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_6_tile_v_1_MPORT_11_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_6_tile_v_1_MPORT_11_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_6_tile_v_0_MPORT_11_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_6_tile_v_0_MPORT_11_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_6_tile_v_0_MPORT_11_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_1_MPORT_156_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_1_MPORT_156_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_1_MPORT_156_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_0_MPORT_156_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_0_MPORT_156_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_0_MPORT_156_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_6_tile_v_3_MPORT_12_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_6_tile_v_3_MPORT_12_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_6_tile_v_3_MPORT_12_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_6_tile_v_2_MPORT_12_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_6_tile_v_2_MPORT_12_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_6_tile_v_2_MPORT_12_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_6_tile_v_1_MPORT_12_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_6_tile_v_1_MPORT_12_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_6_tile_v_1_MPORT_12_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_6_tile_v_0_MPORT_12_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_6_tile_v_0_MPORT_12_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_6_tile_v_0_MPORT_12_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_6_tile_v_3_MPORT_12_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_6_tile_v_3_MPORT_12_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_6_tile_v_3_MPORT_12_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_6_tile_v_2_MPORT_12_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_6_tile_v_2_MPORT_12_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_6_tile_v_2_MPORT_12_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_6_tile_v_1_MPORT_12_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_6_tile_v_1_MPORT_12_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_6_tile_v_1_MPORT_12_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_6_tile_v_0_MPORT_12_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_6_tile_v_0_MPORT_12_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_6_tile_v_0_MPORT_12_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_3_MPORT_52_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_3_MPORT_52_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_3_MPORT_52_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_2_MPORT_52_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_2_MPORT_52_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_2_MPORT_52_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_1_MPORT_157_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_1_MPORT_157_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_1_MPORT_157_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_0_MPORT_157_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_0_MPORT_157_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_0_MPORT_157_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_6_tile_v_3_MPORT_13_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_6_tile_v_3_MPORT_13_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_6_tile_v_3_MPORT_13_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_6_tile_v_2_MPORT_13_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_6_tile_v_2_MPORT_13_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_6_tile_v_2_MPORT_13_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_6_tile_v_1_MPORT_13_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_6_tile_v_1_MPORT_13_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_6_tile_v_1_MPORT_13_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_6_tile_v_0_MPORT_13_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_6_tile_v_0_MPORT_13_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_6_tile_v_0_MPORT_13_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_6_tile_v_3_MPORT_13_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_6_tile_v_3_MPORT_13_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_6_tile_v_3_MPORT_13_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_6_tile_v_2_MPORT_13_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_6_tile_v_2_MPORT_13_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_6_tile_v_2_MPORT_13_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_6_tile_v_1_MPORT_13_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_6_tile_v_1_MPORT_13_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_6_tile_v_1_MPORT_13_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_6_tile_v_0_MPORT_13_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_6_tile_v_0_MPORT_13_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_6_tile_v_0_MPORT_13_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_1_MPORT_158_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_1_MPORT_158_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_1_MPORT_158_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_0_MPORT_158_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_0_MPORT_158_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_0_MPORT_158_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_6_tile_v_3_MPORT_14_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_6_tile_v_3_MPORT_14_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_6_tile_v_3_MPORT_14_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_6_tile_v_2_MPORT_14_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_6_tile_v_2_MPORT_14_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_6_tile_v_2_MPORT_14_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_6_tile_v_1_MPORT_14_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_6_tile_v_1_MPORT_14_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_6_tile_v_1_MPORT_14_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_6_tile_v_0_MPORT_14_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_6_tile_v_0_MPORT_14_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_6_tile_v_0_MPORT_14_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_6_tile_v_3_MPORT_14_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_6_tile_v_3_MPORT_14_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_6_tile_v_3_MPORT_14_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_6_tile_v_2_MPORT_14_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_6_tile_v_2_MPORT_14_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_6_tile_v_2_MPORT_14_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_6_tile_v_1_MPORT_14_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_6_tile_v_1_MPORT_14_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_6_tile_v_1_MPORT_14_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_6_tile_v_0_MPORT_14_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_6_tile_v_0_MPORT_14_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_6_tile_v_0_MPORT_14_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_3_MPORT_53_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_3_MPORT_53_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_3_MPORT_53_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_2_MPORT_53_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_2_MPORT_53_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_2_MPORT_53_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_1_MPORT_159_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_1_MPORT_159_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_1_MPORT_159_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_0_MPORT_159_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_0_MPORT_159_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_0_MPORT_159_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_6_tile_v_3_MPORT_15_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_6_tile_v_3_MPORT_15_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_6_tile_v_3_MPORT_15_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_6_tile_v_2_MPORT_15_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_6_tile_v_2_MPORT_15_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_6_tile_v_2_MPORT_15_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_6_tile_v_1_MPORT_15_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_6_tile_v_1_MPORT_15_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_6_tile_v_1_MPORT_15_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_6_tile_v_0_MPORT_15_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_6_tile_v_0_MPORT_15_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_6_tile_v_0_MPORT_15_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_6_tile_v_3_MPORT_15_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_6_tile_v_3_MPORT_15_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_6_tile_v_3_MPORT_15_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_6_tile_v_2_MPORT_15_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_6_tile_v_2_MPORT_15_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_6_tile_v_2_MPORT_15_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_6_tile_v_1_MPORT_15_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_6_tile_v_1_MPORT_15_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_6_tile_v_1_MPORT_15_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_6_tile_v_0_MPORT_15_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_6_tile_v_0_MPORT_15_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_6_tile_v_0_MPORT_15_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_1_MPORT_160_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_1_MPORT_160_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_1_MPORT_160_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_0_MPORT_160_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_0_MPORT_160_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_0_MPORT_160_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_6_tile_v_3_MPORT_16_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_6_tile_v_3_MPORT_16_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_6_tile_v_3_MPORT_16_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_6_tile_v_2_MPORT_16_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_6_tile_v_2_MPORT_16_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_6_tile_v_2_MPORT_16_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_6_tile_v_1_MPORT_16_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_6_tile_v_1_MPORT_16_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_6_tile_v_1_MPORT_16_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_6_tile_v_0_MPORT_16_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_6_tile_v_0_MPORT_16_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_6_tile_v_0_MPORT_16_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_6_tile_v_3_MPORT_16_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_6_tile_v_3_MPORT_16_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_6_tile_v_3_MPORT_16_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_6_tile_v_2_MPORT_16_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_6_tile_v_2_MPORT_16_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_6_tile_v_2_MPORT_16_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_6_tile_v_1_MPORT_16_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_6_tile_v_1_MPORT_16_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_6_tile_v_1_MPORT_16_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_6_tile_v_0_MPORT_16_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_6_tile_v_0_MPORT_16_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_6_tile_v_0_MPORT_16_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_1_MPORT_161_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_1_MPORT_161_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_1_MPORT_161_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_0_MPORT_161_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_0_MPORT_161_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_0_MPORT_161_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_6_tile_v_3_MPORT_17_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_6_tile_v_3_MPORT_17_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_6_tile_v_3_MPORT_17_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_6_tile_v_2_MPORT_17_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_6_tile_v_2_MPORT_17_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_6_tile_v_2_MPORT_17_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_6_tile_v_1_MPORT_17_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_6_tile_v_1_MPORT_17_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_6_tile_v_1_MPORT_17_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_6_tile_v_0_MPORT_17_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_6_tile_v_0_MPORT_17_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_6_tile_v_0_MPORT_17_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_6_tile_v_3_MPORT_17_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_6_tile_v_3_MPORT_17_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_6_tile_v_3_MPORT_17_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_6_tile_v_2_MPORT_17_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_6_tile_v_2_MPORT_17_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_6_tile_v_2_MPORT_17_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_6_tile_v_1_MPORT_17_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_6_tile_v_1_MPORT_17_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_6_tile_v_1_MPORT_17_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_6_tile_v_0_MPORT_17_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_6_tile_v_0_MPORT_17_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_6_tile_v_0_MPORT_17_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_1_MPORT_162_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_1_MPORT_162_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_1_MPORT_162_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_0_MPORT_162_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_0_MPORT_162_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_0_MPORT_162_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_6_tile_v_3_MPORT_18_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_6_tile_v_3_MPORT_18_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_6_tile_v_3_MPORT_18_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_6_tile_v_2_MPORT_18_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_6_tile_v_2_MPORT_18_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_6_tile_v_2_MPORT_18_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_6_tile_v_1_MPORT_18_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_6_tile_v_1_MPORT_18_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_6_tile_v_1_MPORT_18_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_6_tile_v_0_MPORT_18_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_6_tile_v_0_MPORT_18_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_6_tile_v_0_MPORT_18_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_6_tile_v_3_MPORT_18_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_6_tile_v_3_MPORT_18_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_6_tile_v_3_MPORT_18_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_6_tile_v_2_MPORT_18_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_6_tile_v_2_MPORT_18_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_6_tile_v_2_MPORT_18_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_6_tile_v_1_MPORT_18_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_6_tile_v_1_MPORT_18_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_6_tile_v_1_MPORT_18_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_6_tile_v_0_MPORT_18_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_6_tile_v_0_MPORT_18_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_6_tile_v_0_MPORT_18_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_3_MPORT_54_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_3_MPORT_54_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_3_MPORT_54_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_2_MPORT_54_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_2_MPORT_54_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_2_MPORT_54_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_1_MPORT_163_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_1_MPORT_163_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_1_MPORT_163_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_0_MPORT_163_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_0_MPORT_163_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_0_MPORT_163_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_6_tile_v_3_MPORT_19_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_6_tile_v_3_MPORT_19_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_6_tile_v_3_MPORT_19_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_6_tile_v_2_MPORT_19_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_6_tile_v_2_MPORT_19_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_6_tile_v_2_MPORT_19_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_6_tile_v_1_MPORT_19_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_6_tile_v_1_MPORT_19_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_6_tile_v_1_MPORT_19_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_6_tile_v_0_MPORT_19_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_6_tile_v_0_MPORT_19_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_6_tile_v_0_MPORT_19_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_6_tile_v_3_MPORT_19_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_6_tile_v_3_MPORT_19_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_6_tile_v_3_MPORT_19_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_6_tile_v_2_MPORT_19_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_6_tile_v_2_MPORT_19_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_6_tile_v_2_MPORT_19_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_6_tile_v_1_MPORT_19_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_6_tile_v_1_MPORT_19_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_6_tile_v_1_MPORT_19_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_6_tile_v_0_MPORT_19_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_6_tile_v_0_MPORT_19_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_6_tile_v_0_MPORT_19_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_1_MPORT_164_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_1_MPORT_164_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_1_MPORT_164_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_0_MPORT_164_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_0_MPORT_164_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_0_MPORT_164_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_6_tile_v_3_MPORT_20_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_6_tile_v_3_MPORT_20_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_6_tile_v_3_MPORT_20_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_6_tile_v_2_MPORT_20_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_6_tile_v_2_MPORT_20_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_6_tile_v_2_MPORT_20_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_6_tile_v_1_MPORT_20_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_6_tile_v_1_MPORT_20_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_6_tile_v_1_MPORT_20_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_6_tile_v_0_MPORT_20_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_6_tile_v_0_MPORT_20_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_6_tile_v_0_MPORT_20_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_6_tile_v_3_MPORT_20_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_6_tile_v_3_MPORT_20_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_6_tile_v_3_MPORT_20_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_6_tile_v_2_MPORT_20_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_6_tile_v_2_MPORT_20_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_6_tile_v_2_MPORT_20_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_6_tile_v_1_MPORT_20_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_6_tile_v_1_MPORT_20_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_6_tile_v_1_MPORT_20_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_6_tile_v_0_MPORT_20_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_6_tile_v_0_MPORT_20_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_6_tile_v_0_MPORT_20_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_3_MPORT_55_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_3_MPORT_55_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_3_MPORT_55_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_2_MPORT_55_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_2_MPORT_55_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_2_MPORT_55_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_1_MPORT_165_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_1_MPORT_165_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_1_MPORT_165_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_0_MPORT_165_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_0_MPORT_165_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_0_MPORT_165_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_6_tile_v_3_MPORT_21_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_6_tile_v_3_MPORT_21_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_6_tile_v_3_MPORT_21_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_6_tile_v_2_MPORT_21_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_6_tile_v_2_MPORT_21_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_6_tile_v_2_MPORT_21_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_6_tile_v_1_MPORT_21_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_6_tile_v_1_MPORT_21_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_6_tile_v_1_MPORT_21_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_6_tile_v_0_MPORT_21_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_6_tile_v_0_MPORT_21_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_6_tile_v_0_MPORT_21_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_6_tile_v_3_MPORT_21_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_6_tile_v_3_MPORT_21_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_6_tile_v_3_MPORT_21_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_6_tile_v_2_MPORT_21_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_6_tile_v_2_MPORT_21_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_6_tile_v_2_MPORT_21_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_6_tile_v_1_MPORT_21_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_6_tile_v_1_MPORT_21_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_6_tile_v_1_MPORT_21_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_6_tile_v_0_MPORT_21_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_6_tile_v_0_MPORT_21_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_6_tile_v_0_MPORT_21_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_1_MPORT_166_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_1_MPORT_166_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_1_MPORT_166_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_0_MPORT_166_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_0_MPORT_166_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_0_MPORT_166_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_6_tile_v_3_MPORT_22_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_6_tile_v_3_MPORT_22_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_6_tile_v_3_MPORT_22_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_6_tile_v_2_MPORT_22_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_6_tile_v_2_MPORT_22_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_6_tile_v_2_MPORT_22_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_6_tile_v_1_MPORT_22_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_6_tile_v_1_MPORT_22_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_6_tile_v_1_MPORT_22_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_6_tile_v_0_MPORT_22_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_6_tile_v_0_MPORT_22_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_6_tile_v_0_MPORT_22_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_6_tile_v_3_MPORT_22_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_6_tile_v_3_MPORT_22_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_6_tile_v_3_MPORT_22_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_6_tile_v_2_MPORT_22_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_6_tile_v_2_MPORT_22_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_6_tile_v_2_MPORT_22_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_6_tile_v_1_MPORT_22_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_6_tile_v_1_MPORT_22_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_6_tile_v_1_MPORT_22_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_6_tile_v_0_MPORT_22_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_6_tile_v_0_MPORT_22_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_6_tile_v_0_MPORT_22_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_1_MPORT_167_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_1_MPORT_167_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_1_MPORT_167_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_0_MPORT_167_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_0_MPORT_167_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_0_MPORT_167_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_6_tile_v_3_MPORT_23_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_6_tile_v_3_MPORT_23_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_6_tile_v_3_MPORT_23_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_6_tile_v_2_MPORT_23_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_6_tile_v_2_MPORT_23_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_6_tile_v_2_MPORT_23_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_6_tile_v_1_MPORT_23_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_6_tile_v_1_MPORT_23_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_6_tile_v_1_MPORT_23_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_6_tile_v_0_MPORT_23_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_6_tile_v_0_MPORT_23_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_6_tile_v_0_MPORT_23_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_6_tile_v_3_MPORT_23_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_6_tile_v_3_MPORT_23_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_6_tile_v_3_MPORT_23_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_6_tile_v_2_MPORT_23_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_6_tile_v_2_MPORT_23_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_6_tile_v_2_MPORT_23_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_6_tile_v_1_MPORT_23_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_6_tile_v_1_MPORT_23_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_6_tile_v_1_MPORT_23_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_6_tile_v_0_MPORT_23_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_6_tile_v_0_MPORT_23_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_6_tile_v_0_MPORT_23_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_1_MPORT_168_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_1_MPORT_168_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_1_MPORT_168_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_0_MPORT_168_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_0_MPORT_168_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_0_MPORT_168_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_7_tile_v_3_MPORT_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_7_tile_v_3_MPORT_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_7_tile_v_3_MPORT_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_7_tile_v_2_MPORT_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_7_tile_v_2_MPORT_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_7_tile_v_2_MPORT_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_7_tile_v_1_MPORT_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_7_tile_v_1_MPORT_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_7_tile_v_1_MPORT_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_7_tile_v_0_MPORT_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_7_tile_v_0_MPORT_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_7_tile_v_0_MPORT_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_7_tile_v_3_MPORT_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_7_tile_v_3_MPORT_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_7_tile_v_3_MPORT_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_7_tile_v_2_MPORT_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_7_tile_v_2_MPORT_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_7_tile_v_2_MPORT_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_7_tile_v_1_MPORT_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_7_tile_v_1_MPORT_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_7_tile_v_1_MPORT_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_7_tile_v_0_MPORT_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_7_tile_v_0_MPORT_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_7_tile_v_0_MPORT_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_3_MPORT_56_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_3_MPORT_56_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_3_MPORT_56_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_2_MPORT_56_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_2_MPORT_56_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_2_MPORT_56_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_1_MPORT_169_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_1_MPORT_169_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_1_MPORT_169_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_0_MPORT_169_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_0_MPORT_169_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_0_MPORT_169_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_7_tile_v_3_MPORT_1_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_7_tile_v_3_MPORT_1_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_7_tile_v_3_MPORT_1_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_7_tile_v_2_MPORT_1_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_7_tile_v_2_MPORT_1_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_7_tile_v_2_MPORT_1_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_7_tile_v_1_MPORT_1_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_7_tile_v_1_MPORT_1_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_7_tile_v_1_MPORT_1_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_7_tile_v_0_MPORT_1_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_7_tile_v_0_MPORT_1_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_7_tile_v_0_MPORT_1_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_7_tile_v_3_MPORT_1_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_7_tile_v_3_MPORT_1_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_7_tile_v_3_MPORT_1_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_7_tile_v_2_MPORT_1_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_7_tile_v_2_MPORT_1_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_7_tile_v_2_MPORT_1_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_7_tile_v_1_MPORT_1_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_7_tile_v_1_MPORT_1_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_7_tile_v_1_MPORT_1_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_7_tile_v_0_MPORT_1_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_7_tile_v_0_MPORT_1_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_7_tile_v_0_MPORT_1_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_1_MPORT_170_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_1_MPORT_170_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_1_MPORT_170_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_0_MPORT_170_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_0_MPORT_170_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_0_MPORT_170_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_7_tile_v_3_MPORT_2_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_7_tile_v_3_MPORT_2_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_7_tile_v_3_MPORT_2_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_7_tile_v_2_MPORT_2_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_7_tile_v_2_MPORT_2_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_7_tile_v_2_MPORT_2_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_7_tile_v_1_MPORT_2_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_7_tile_v_1_MPORT_2_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_7_tile_v_1_MPORT_2_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_7_tile_v_0_MPORT_2_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_7_tile_v_0_MPORT_2_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_7_tile_v_0_MPORT_2_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_7_tile_v_3_MPORT_2_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_7_tile_v_3_MPORT_2_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_7_tile_v_3_MPORT_2_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_7_tile_v_2_MPORT_2_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_7_tile_v_2_MPORT_2_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_7_tile_v_2_MPORT_2_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_7_tile_v_1_MPORT_2_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_7_tile_v_1_MPORT_2_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_7_tile_v_1_MPORT_2_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_7_tile_v_0_MPORT_2_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_7_tile_v_0_MPORT_2_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_7_tile_v_0_MPORT_2_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_3_MPORT_57_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_3_MPORT_57_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_3_MPORT_57_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_2_MPORT_57_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_2_MPORT_57_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_2_MPORT_57_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_1_MPORT_171_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_1_MPORT_171_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_1_MPORT_171_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_0_MPORT_171_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_0_MPORT_171_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_0_MPORT_171_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_7_tile_v_3_MPORT_3_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_7_tile_v_3_MPORT_3_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_7_tile_v_3_MPORT_3_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_7_tile_v_2_MPORT_3_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_7_tile_v_2_MPORT_3_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_7_tile_v_2_MPORT_3_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_7_tile_v_1_MPORT_3_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_7_tile_v_1_MPORT_3_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_7_tile_v_1_MPORT_3_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_7_tile_v_0_MPORT_3_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_7_tile_v_0_MPORT_3_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_7_tile_v_0_MPORT_3_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_7_tile_v_3_MPORT_3_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_7_tile_v_3_MPORT_3_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_7_tile_v_3_MPORT_3_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_7_tile_v_2_MPORT_3_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_7_tile_v_2_MPORT_3_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_7_tile_v_2_MPORT_3_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_7_tile_v_1_MPORT_3_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_7_tile_v_1_MPORT_3_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_7_tile_v_1_MPORT_3_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_7_tile_v_0_MPORT_3_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_7_tile_v_0_MPORT_3_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_7_tile_v_0_MPORT_3_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_1_MPORT_172_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_1_MPORT_172_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_1_MPORT_172_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_0_MPORT_172_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_0_MPORT_172_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_0_MPORT_172_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_7_tile_v_3_MPORT_4_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_7_tile_v_3_MPORT_4_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_7_tile_v_3_MPORT_4_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_7_tile_v_2_MPORT_4_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_7_tile_v_2_MPORT_4_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_7_tile_v_2_MPORT_4_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_7_tile_v_1_MPORT_4_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_7_tile_v_1_MPORT_4_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_7_tile_v_1_MPORT_4_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_7_tile_v_0_MPORT_4_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_7_tile_v_0_MPORT_4_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_7_tile_v_0_MPORT_4_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_7_tile_v_3_MPORT_4_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_7_tile_v_3_MPORT_4_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_7_tile_v_3_MPORT_4_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_7_tile_v_2_MPORT_4_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_7_tile_v_2_MPORT_4_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_7_tile_v_2_MPORT_4_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_7_tile_v_1_MPORT_4_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_7_tile_v_1_MPORT_4_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_7_tile_v_1_MPORT_4_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_7_tile_v_0_MPORT_4_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_7_tile_v_0_MPORT_4_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_7_tile_v_0_MPORT_4_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_1_MPORT_173_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_1_MPORT_173_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_1_MPORT_173_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_0_MPORT_173_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_0_MPORT_173_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_0_MPORT_173_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_7_tile_v_3_MPORT_5_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_7_tile_v_3_MPORT_5_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_7_tile_v_3_MPORT_5_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_7_tile_v_2_MPORT_5_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_7_tile_v_2_MPORT_5_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_7_tile_v_2_MPORT_5_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_7_tile_v_1_MPORT_5_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_7_tile_v_1_MPORT_5_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_7_tile_v_1_MPORT_5_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_7_tile_v_0_MPORT_5_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_7_tile_v_0_MPORT_5_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_7_tile_v_0_MPORT_5_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_7_tile_v_3_MPORT_5_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_7_tile_v_3_MPORT_5_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_7_tile_v_3_MPORT_5_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_7_tile_v_2_MPORT_5_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_7_tile_v_2_MPORT_5_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_7_tile_v_2_MPORT_5_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_7_tile_v_1_MPORT_5_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_7_tile_v_1_MPORT_5_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_7_tile_v_1_MPORT_5_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_7_tile_v_0_MPORT_5_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_7_tile_v_0_MPORT_5_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_7_tile_v_0_MPORT_5_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_1_MPORT_174_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_1_MPORT_174_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_1_MPORT_174_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_0_MPORT_174_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_0_MPORT_174_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_0_MPORT_174_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_7_tile_v_3_MPORT_6_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_7_tile_v_3_MPORT_6_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_7_tile_v_3_MPORT_6_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_7_tile_v_2_MPORT_6_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_7_tile_v_2_MPORT_6_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_7_tile_v_2_MPORT_6_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_7_tile_v_1_MPORT_6_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_7_tile_v_1_MPORT_6_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_7_tile_v_1_MPORT_6_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_7_tile_v_0_MPORT_6_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_7_tile_v_0_MPORT_6_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_7_tile_v_0_MPORT_6_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_7_tile_v_3_MPORT_6_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_7_tile_v_3_MPORT_6_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_7_tile_v_3_MPORT_6_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_7_tile_v_2_MPORT_6_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_7_tile_v_2_MPORT_6_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_7_tile_v_2_MPORT_6_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_7_tile_v_1_MPORT_6_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_7_tile_v_1_MPORT_6_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_7_tile_v_1_MPORT_6_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_7_tile_v_0_MPORT_6_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_7_tile_v_0_MPORT_6_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_7_tile_v_0_MPORT_6_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_3_MPORT_58_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_3_MPORT_58_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_3_MPORT_58_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_2_MPORT_58_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_2_MPORT_58_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_2_MPORT_58_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_1_MPORT_175_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_1_MPORT_175_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_1_MPORT_175_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_0_MPORT_175_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_0_MPORT_175_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_0_MPORT_175_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_7_tile_v_3_MPORT_7_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_7_tile_v_3_MPORT_7_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_7_tile_v_3_MPORT_7_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_7_tile_v_2_MPORT_7_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_7_tile_v_2_MPORT_7_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_7_tile_v_2_MPORT_7_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_7_tile_v_1_MPORT_7_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_7_tile_v_1_MPORT_7_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_7_tile_v_1_MPORT_7_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_7_tile_v_0_MPORT_7_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_7_tile_v_0_MPORT_7_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_7_tile_v_0_MPORT_7_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_7_tile_v_3_MPORT_7_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_7_tile_v_3_MPORT_7_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_7_tile_v_3_MPORT_7_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_7_tile_v_2_MPORT_7_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_7_tile_v_2_MPORT_7_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_7_tile_v_2_MPORT_7_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_7_tile_v_1_MPORT_7_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_7_tile_v_1_MPORT_7_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_7_tile_v_1_MPORT_7_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_7_tile_v_0_MPORT_7_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_7_tile_v_0_MPORT_7_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_7_tile_v_0_MPORT_7_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_1_MPORT_176_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_1_MPORT_176_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_1_MPORT_176_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_0_MPORT_176_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_0_MPORT_176_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_0_MPORT_176_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_7_tile_v_3_MPORT_8_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_7_tile_v_3_MPORT_8_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_7_tile_v_3_MPORT_8_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_7_tile_v_2_MPORT_8_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_7_tile_v_2_MPORT_8_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_7_tile_v_2_MPORT_8_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_7_tile_v_1_MPORT_8_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_7_tile_v_1_MPORT_8_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_7_tile_v_1_MPORT_8_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_7_tile_v_0_MPORT_8_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_7_tile_v_0_MPORT_8_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_7_tile_v_0_MPORT_8_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_7_tile_v_3_MPORT_8_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_7_tile_v_3_MPORT_8_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_7_tile_v_3_MPORT_8_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_7_tile_v_2_MPORT_8_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_7_tile_v_2_MPORT_8_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_7_tile_v_2_MPORT_8_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_7_tile_v_1_MPORT_8_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_7_tile_v_1_MPORT_8_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_7_tile_v_1_MPORT_8_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_7_tile_v_0_MPORT_8_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_7_tile_v_0_MPORT_8_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_7_tile_v_0_MPORT_8_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_3_MPORT_59_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_3_MPORT_59_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_3_MPORT_59_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_2_MPORT_59_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_2_MPORT_59_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_2_MPORT_59_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_1_MPORT_177_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_1_MPORT_177_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_1_MPORT_177_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_0_MPORT_177_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_0_MPORT_177_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_0_MPORT_177_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_7_tile_v_3_MPORT_9_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_7_tile_v_3_MPORT_9_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_7_tile_v_3_MPORT_9_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_7_tile_v_2_MPORT_9_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_7_tile_v_2_MPORT_9_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_7_tile_v_2_MPORT_9_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_7_tile_v_1_MPORT_9_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_7_tile_v_1_MPORT_9_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_7_tile_v_1_MPORT_9_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_7_tile_v_0_MPORT_9_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_7_tile_v_0_MPORT_9_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_7_tile_v_0_MPORT_9_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_7_tile_v_3_MPORT_9_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_7_tile_v_3_MPORT_9_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_7_tile_v_3_MPORT_9_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_7_tile_v_2_MPORT_9_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_7_tile_v_2_MPORT_9_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_7_tile_v_2_MPORT_9_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_7_tile_v_1_MPORT_9_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_7_tile_v_1_MPORT_9_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_7_tile_v_1_MPORT_9_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_7_tile_v_0_MPORT_9_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_7_tile_v_0_MPORT_9_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_7_tile_v_0_MPORT_9_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_1_MPORT_178_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_1_MPORT_178_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_1_MPORT_178_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_0_MPORT_178_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_0_MPORT_178_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_0_MPORT_178_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_7_tile_v_3_MPORT_10_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_7_tile_v_3_MPORT_10_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_7_tile_v_3_MPORT_10_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_7_tile_v_2_MPORT_10_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_7_tile_v_2_MPORT_10_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_7_tile_v_2_MPORT_10_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_7_tile_v_1_MPORT_10_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_7_tile_v_1_MPORT_10_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_7_tile_v_1_MPORT_10_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_7_tile_v_0_MPORT_10_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_7_tile_v_0_MPORT_10_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_7_tile_v_0_MPORT_10_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_7_tile_v_3_MPORT_10_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_7_tile_v_3_MPORT_10_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_7_tile_v_3_MPORT_10_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_7_tile_v_2_MPORT_10_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_7_tile_v_2_MPORT_10_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_7_tile_v_2_MPORT_10_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_7_tile_v_1_MPORT_10_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_7_tile_v_1_MPORT_10_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_7_tile_v_1_MPORT_10_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_7_tile_v_0_MPORT_10_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_7_tile_v_0_MPORT_10_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_7_tile_v_0_MPORT_10_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_1_MPORT_179_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_1_MPORT_179_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_1_MPORT_179_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_0_MPORT_179_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_0_MPORT_179_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_0_MPORT_179_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_7_tile_v_3_MPORT_11_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_7_tile_v_3_MPORT_11_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_7_tile_v_3_MPORT_11_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_7_tile_v_2_MPORT_11_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_7_tile_v_2_MPORT_11_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_7_tile_v_2_MPORT_11_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_7_tile_v_1_MPORT_11_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_7_tile_v_1_MPORT_11_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_7_tile_v_1_MPORT_11_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_7_tile_v_0_MPORT_11_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_7_tile_v_0_MPORT_11_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_7_tile_v_0_MPORT_11_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_7_tile_v_3_MPORT_11_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_7_tile_v_3_MPORT_11_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_7_tile_v_3_MPORT_11_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_7_tile_v_2_MPORT_11_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_7_tile_v_2_MPORT_11_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_7_tile_v_2_MPORT_11_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_7_tile_v_1_MPORT_11_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_7_tile_v_1_MPORT_11_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_7_tile_v_1_MPORT_11_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_7_tile_v_0_MPORT_11_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_7_tile_v_0_MPORT_11_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_7_tile_v_0_MPORT_11_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_1_MPORT_180_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_1_MPORT_180_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_1_MPORT_180_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_0_MPORT_180_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_0_MPORT_180_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_0_MPORT_180_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_7_tile_v_3_MPORT_12_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_7_tile_v_3_MPORT_12_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_7_tile_v_3_MPORT_12_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_7_tile_v_2_MPORT_12_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_7_tile_v_2_MPORT_12_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_7_tile_v_2_MPORT_12_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_7_tile_v_1_MPORT_12_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_7_tile_v_1_MPORT_12_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_7_tile_v_1_MPORT_12_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_7_tile_v_0_MPORT_12_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_7_tile_v_0_MPORT_12_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_7_tile_v_0_MPORT_12_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_7_tile_v_3_MPORT_12_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_7_tile_v_3_MPORT_12_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_7_tile_v_3_MPORT_12_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_7_tile_v_2_MPORT_12_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_7_tile_v_2_MPORT_12_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_7_tile_v_2_MPORT_12_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_7_tile_v_1_MPORT_12_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_7_tile_v_1_MPORT_12_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_7_tile_v_1_MPORT_12_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_7_tile_v_0_MPORT_12_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_7_tile_v_0_MPORT_12_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_7_tile_v_0_MPORT_12_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_3_MPORT_60_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_3_MPORT_60_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_3_MPORT_60_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_2_MPORT_60_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_2_MPORT_60_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_2_MPORT_60_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_1_MPORT_181_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_1_MPORT_181_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_1_MPORT_181_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_0_MPORT_181_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_0_MPORT_181_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_0_MPORT_181_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_7_tile_v_3_MPORT_13_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_7_tile_v_3_MPORT_13_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_7_tile_v_3_MPORT_13_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_7_tile_v_2_MPORT_13_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_7_tile_v_2_MPORT_13_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_7_tile_v_2_MPORT_13_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_7_tile_v_1_MPORT_13_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_7_tile_v_1_MPORT_13_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_7_tile_v_1_MPORT_13_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_7_tile_v_0_MPORT_13_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_7_tile_v_0_MPORT_13_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_7_tile_v_0_MPORT_13_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_7_tile_v_3_MPORT_13_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_7_tile_v_3_MPORT_13_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_7_tile_v_3_MPORT_13_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_7_tile_v_2_MPORT_13_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_7_tile_v_2_MPORT_13_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_7_tile_v_2_MPORT_13_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_7_tile_v_1_MPORT_13_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_7_tile_v_1_MPORT_13_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_7_tile_v_1_MPORT_13_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_7_tile_v_0_MPORT_13_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_7_tile_v_0_MPORT_13_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_7_tile_v_0_MPORT_13_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_1_MPORT_182_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_1_MPORT_182_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_1_MPORT_182_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_0_MPORT_182_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_0_MPORT_182_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_0_MPORT_182_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_7_tile_v_3_MPORT_14_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_7_tile_v_3_MPORT_14_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_7_tile_v_3_MPORT_14_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_7_tile_v_2_MPORT_14_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_7_tile_v_2_MPORT_14_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_7_tile_v_2_MPORT_14_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_7_tile_v_1_MPORT_14_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_7_tile_v_1_MPORT_14_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_7_tile_v_1_MPORT_14_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_7_tile_v_0_MPORT_14_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_7_tile_v_0_MPORT_14_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_7_tile_v_0_MPORT_14_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_7_tile_v_3_MPORT_14_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_7_tile_v_3_MPORT_14_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_7_tile_v_3_MPORT_14_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_7_tile_v_2_MPORT_14_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_7_tile_v_2_MPORT_14_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_7_tile_v_2_MPORT_14_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_7_tile_v_1_MPORT_14_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_7_tile_v_1_MPORT_14_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_7_tile_v_1_MPORT_14_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_7_tile_v_0_MPORT_14_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_7_tile_v_0_MPORT_14_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_7_tile_v_0_MPORT_14_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_3_MPORT_61_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_3_MPORT_61_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_3_MPORT_61_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_2_MPORT_61_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_2_MPORT_61_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_2_MPORT_61_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_1_MPORT_183_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_1_MPORT_183_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_1_MPORT_183_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_0_MPORT_183_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_0_MPORT_183_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_0_MPORT_183_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_7_tile_v_3_MPORT_15_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_7_tile_v_3_MPORT_15_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_7_tile_v_3_MPORT_15_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_7_tile_v_2_MPORT_15_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_7_tile_v_2_MPORT_15_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_7_tile_v_2_MPORT_15_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_7_tile_v_1_MPORT_15_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_7_tile_v_1_MPORT_15_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_7_tile_v_1_MPORT_15_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_7_tile_v_0_MPORT_15_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_7_tile_v_0_MPORT_15_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_7_tile_v_0_MPORT_15_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_7_tile_v_3_MPORT_15_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_7_tile_v_3_MPORT_15_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_7_tile_v_3_MPORT_15_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_7_tile_v_2_MPORT_15_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_7_tile_v_2_MPORT_15_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_7_tile_v_2_MPORT_15_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_7_tile_v_1_MPORT_15_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_7_tile_v_1_MPORT_15_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_7_tile_v_1_MPORT_15_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_7_tile_v_0_MPORT_15_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_7_tile_v_0_MPORT_15_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_7_tile_v_0_MPORT_15_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_1_MPORT_184_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_1_MPORT_184_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_1_MPORT_184_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_0_MPORT_184_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_0_MPORT_184_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_0_MPORT_184_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_7_tile_v_3_MPORT_16_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_7_tile_v_3_MPORT_16_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_7_tile_v_3_MPORT_16_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_7_tile_v_2_MPORT_16_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_7_tile_v_2_MPORT_16_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_7_tile_v_2_MPORT_16_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_7_tile_v_1_MPORT_16_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_7_tile_v_1_MPORT_16_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_7_tile_v_1_MPORT_16_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_7_tile_v_0_MPORT_16_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_7_tile_v_0_MPORT_16_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_7_tile_v_0_MPORT_16_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_7_tile_v_3_MPORT_16_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_7_tile_v_3_MPORT_16_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_7_tile_v_3_MPORT_16_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_7_tile_v_2_MPORT_16_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_7_tile_v_2_MPORT_16_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_7_tile_v_2_MPORT_16_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_7_tile_v_1_MPORT_16_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_7_tile_v_1_MPORT_16_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_7_tile_v_1_MPORT_16_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_7_tile_v_0_MPORT_16_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_7_tile_v_0_MPORT_16_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_7_tile_v_0_MPORT_16_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_1_MPORT_185_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_1_MPORT_185_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_1_MPORT_185_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_0_MPORT_185_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_0_MPORT_185_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_0_MPORT_185_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_7_tile_v_3_MPORT_17_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_7_tile_v_3_MPORT_17_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_7_tile_v_3_MPORT_17_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_7_tile_v_2_MPORT_17_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_7_tile_v_2_MPORT_17_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_7_tile_v_2_MPORT_17_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_7_tile_v_1_MPORT_17_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_7_tile_v_1_MPORT_17_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_7_tile_v_1_MPORT_17_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_7_tile_v_0_MPORT_17_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_7_tile_v_0_MPORT_17_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_7_tile_v_0_MPORT_17_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_7_tile_v_3_MPORT_17_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_7_tile_v_3_MPORT_17_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_7_tile_v_3_MPORT_17_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_7_tile_v_2_MPORT_17_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_7_tile_v_2_MPORT_17_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_7_tile_v_2_MPORT_17_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_7_tile_v_1_MPORT_17_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_7_tile_v_1_MPORT_17_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_7_tile_v_1_MPORT_17_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_7_tile_v_0_MPORT_17_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_7_tile_v_0_MPORT_17_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_7_tile_v_0_MPORT_17_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_1_MPORT_186_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_1_MPORT_186_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_1_MPORT_186_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_0_MPORT_186_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_0_MPORT_186_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_0_MPORT_186_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_7_tile_v_3_MPORT_18_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_7_tile_v_3_MPORT_18_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_7_tile_v_3_MPORT_18_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_7_tile_v_2_MPORT_18_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_7_tile_v_2_MPORT_18_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_7_tile_v_2_MPORT_18_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_7_tile_v_1_MPORT_18_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_7_tile_v_1_MPORT_18_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_7_tile_v_1_MPORT_18_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_7_tile_v_0_MPORT_18_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_7_tile_v_0_MPORT_18_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_7_tile_v_0_MPORT_18_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_7_tile_v_3_MPORT_18_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_7_tile_v_3_MPORT_18_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_7_tile_v_3_MPORT_18_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_7_tile_v_2_MPORT_18_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_7_tile_v_2_MPORT_18_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_7_tile_v_2_MPORT_18_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_7_tile_v_1_MPORT_18_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_7_tile_v_1_MPORT_18_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_7_tile_v_1_MPORT_18_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_7_tile_v_0_MPORT_18_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_7_tile_v_0_MPORT_18_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_7_tile_v_0_MPORT_18_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_3_MPORT_62_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_3_MPORT_62_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_3_MPORT_62_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_2_MPORT_62_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_2_MPORT_62_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_2_MPORT_62_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_1_MPORT_187_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_1_MPORT_187_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_1_MPORT_187_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_0_MPORT_187_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_0_MPORT_187_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_0_MPORT_187_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_7_tile_v_3_MPORT_19_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_7_tile_v_3_MPORT_19_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_7_tile_v_3_MPORT_19_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_7_tile_v_2_MPORT_19_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_7_tile_v_2_MPORT_19_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_7_tile_v_2_MPORT_19_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_7_tile_v_1_MPORT_19_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_7_tile_v_1_MPORT_19_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_7_tile_v_1_MPORT_19_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_7_tile_v_0_MPORT_19_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_7_tile_v_0_MPORT_19_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_7_tile_v_0_MPORT_19_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_7_tile_v_3_MPORT_19_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_7_tile_v_3_MPORT_19_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_7_tile_v_3_MPORT_19_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_7_tile_v_2_MPORT_19_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_7_tile_v_2_MPORT_19_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_7_tile_v_2_MPORT_19_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_7_tile_v_1_MPORT_19_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_7_tile_v_1_MPORT_19_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_7_tile_v_1_MPORT_19_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_7_tile_v_0_MPORT_19_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_7_tile_v_0_MPORT_19_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_7_tile_v_0_MPORT_19_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_1_MPORT_188_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_1_MPORT_188_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_1_MPORT_188_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_0_MPORT_188_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_0_MPORT_188_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_0_MPORT_188_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_7_tile_v_3_MPORT_20_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_7_tile_v_3_MPORT_20_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_7_tile_v_3_MPORT_20_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_7_tile_v_2_MPORT_20_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_7_tile_v_2_MPORT_20_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_7_tile_v_2_MPORT_20_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_7_tile_v_1_MPORT_20_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_7_tile_v_1_MPORT_20_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_7_tile_v_1_MPORT_20_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_7_tile_v_0_MPORT_20_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_7_tile_v_0_MPORT_20_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_7_tile_v_0_MPORT_20_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_7_tile_v_3_MPORT_20_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_7_tile_v_3_MPORT_20_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_7_tile_v_3_MPORT_20_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_7_tile_v_2_MPORT_20_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_7_tile_v_2_MPORT_20_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_7_tile_v_2_MPORT_20_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_7_tile_v_1_MPORT_20_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_7_tile_v_1_MPORT_20_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_7_tile_v_1_MPORT_20_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_7_tile_v_0_MPORT_20_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_7_tile_v_0_MPORT_20_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_7_tile_v_0_MPORT_20_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_3_MPORT_63_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_3_MPORT_63_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_3_MPORT_63_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_2_MPORT_63_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_2_MPORT_63_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_2_MPORT_63_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_1_MPORT_189_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_1_MPORT_189_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_1_MPORT_189_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_0_MPORT_189_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_0_MPORT_189_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_0_MPORT_189_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_7_tile_v_3_MPORT_21_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_7_tile_v_3_MPORT_21_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_7_tile_v_3_MPORT_21_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_7_tile_v_2_MPORT_21_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_7_tile_v_2_MPORT_21_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_7_tile_v_2_MPORT_21_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_7_tile_v_1_MPORT_21_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_7_tile_v_1_MPORT_21_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_7_tile_v_1_MPORT_21_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_7_tile_v_0_MPORT_21_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_7_tile_v_0_MPORT_21_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_7_tile_v_0_MPORT_21_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_7_tile_v_3_MPORT_21_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_7_tile_v_3_MPORT_21_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_7_tile_v_3_MPORT_21_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_7_tile_v_2_MPORT_21_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_7_tile_v_2_MPORT_21_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_7_tile_v_2_MPORT_21_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_7_tile_v_1_MPORT_21_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_7_tile_v_1_MPORT_21_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_7_tile_v_1_MPORT_21_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_7_tile_v_0_MPORT_21_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_7_tile_v_0_MPORT_21_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_7_tile_v_0_MPORT_21_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_1_MPORT_190_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_1_MPORT_190_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_1_MPORT_190_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_0_MPORT_190_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_0_MPORT_190_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_0_MPORT_190_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_7_tile_v_3_MPORT_22_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_7_tile_v_3_MPORT_22_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_7_tile_v_3_MPORT_22_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_7_tile_v_2_MPORT_22_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_7_tile_v_2_MPORT_22_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_7_tile_v_2_MPORT_22_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_7_tile_v_1_MPORT_22_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_7_tile_v_1_MPORT_22_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_7_tile_v_1_MPORT_22_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_7_tile_v_0_MPORT_22_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_7_tile_v_0_MPORT_22_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_7_tile_v_0_MPORT_22_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_7_tile_v_3_MPORT_22_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_7_tile_v_3_MPORT_22_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_7_tile_v_3_MPORT_22_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_7_tile_v_2_MPORT_22_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_7_tile_v_2_MPORT_22_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_7_tile_v_2_MPORT_22_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_7_tile_v_1_MPORT_22_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_7_tile_v_1_MPORT_22_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_7_tile_v_1_MPORT_22_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_7_tile_v_0_MPORT_22_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_7_tile_v_0_MPORT_22_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_7_tile_v_0_MPORT_22_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_1_MPORT_191_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_1_MPORT_191_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_1_MPORT_191_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_a_tile_v_0_MPORT_191_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_a_tile_v_0_MPORT_191_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_a_tile_v_0_MPORT_191_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_7_tile_v_3_MPORT_23_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_7_tile_v_3_MPORT_23_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_7_tile_v_3_MPORT_23_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_7_tile_v_2_MPORT_23_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_7_tile_v_2_MPORT_23_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_7_tile_v_2_MPORT_23_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_7_tile_v_1_MPORT_23_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_7_tile_v_1_MPORT_23_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_7_tile_v_1_MPORT_23_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_b_7_tile_v_0_MPORT_23_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_b_7_tile_v_0_MPORT_23_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_b_7_tile_v_0_MPORT_23_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_7_tile_v_3_MPORT_23_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_7_tile_v_3_MPORT_23_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_7_tile_v_3_MPORT_23_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_7_tile_v_2_MPORT_23_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_7_tile_v_2_MPORT_23_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_7_tile_v_2_MPORT_23_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_7_tile_v_1_MPORT_23_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_7_tile_v_1_MPORT_23_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_7_tile_v_1_MPORT_23_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_matrix_c_7_tile_v_0_MPORT_23_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_matrix_c_7_tile_v_0_MPORT_23_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_matrix_c_7_tile_v_0_MPORT_23_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_io_uart_rf_r_data_MPORT_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_io_uart_rf_r_data_MPORT_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_io_uart_rf_r_data_MPORT_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_MPORT_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_MPORT_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_mask; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_MPORT_1_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_MPORT_1_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_1_mask; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_1_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_MPORT_2_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_MPORT_2_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_2_mask; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_2_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_MPORT_3_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_MPORT_3_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_3_mask; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_3_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_MPORT_4_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_MPORT_4_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_4_mask; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_4_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_MPORT_5_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_MPORT_5_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_5_mask; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_5_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_MPORT_6_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_MPORT_6_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_6_mask; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_6_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_MPORT_7_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_MPORT_7_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_7_mask; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_7_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_MPORT_8_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_MPORT_8_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_8_mask; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_8_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_MPORT_9_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_MPORT_9_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_9_mask; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_9_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_MPORT_10_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_MPORT_10_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_10_mask; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_10_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_MPORT_11_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_MPORT_11_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_11_mask; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_11_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_MPORT_12_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_MPORT_12_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_12_mask; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_12_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_MPORT_13_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_MPORT_13_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_13_mask; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_13_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_MPORT_14_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_MPORT_14_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_14_mask; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_14_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_MPORT_15_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_MPORT_15_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_15_mask; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_15_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_MPORT_16_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_MPORT_16_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_16_mask; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_16_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_MPORT_17_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_MPORT_17_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_17_mask; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_17_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_MPORT_18_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_MPORT_18_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_18_mask; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_18_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_MPORT_19_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_MPORT_19_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_19_mask; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_19_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_MPORT_20_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_MPORT_20_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_20_mask; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_20_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_MPORT_21_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_MPORT_21_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_21_mask; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_21_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_MPORT_22_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_MPORT_22_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_22_mask; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_22_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_MPORT_23_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_MPORT_23_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_23_mask; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_23_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_MPORT_24_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_MPORT_24_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_24_mask; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_24_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_MPORT_25_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_MPORT_25_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_25_mask; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_25_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_MPORT_26_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_MPORT_26_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_26_mask; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_26_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_MPORT_27_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_MPORT_27_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_27_mask; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_27_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_MPORT_28_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_MPORT_28_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_28_mask; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_28_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_MPORT_29_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_MPORT_29_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_29_mask; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_29_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_MPORT_30_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_MPORT_30_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_30_mask; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_30_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_MPORT_31_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_MPORT_31_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_31_mask; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_31_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_MPORT_32_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_MPORT_32_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_32_mask; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_32_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_MPORT_33_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_MPORT_33_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_33_mask; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_33_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_MPORT_34_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_MPORT_34_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_34_mask; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_34_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_MPORT_35_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_MPORT_35_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_35_mask; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_35_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_MPORT_36_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_MPORT_36_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_36_mask; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_36_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_MPORT_37_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_MPORT_37_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_37_mask; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_37_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_MPORT_38_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_MPORT_38_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_38_mask; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_38_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_MPORT_39_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_MPORT_39_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_39_mask; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_39_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_MPORT_40_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_MPORT_40_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_40_mask; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_40_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_MPORT_41_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_MPORT_41_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_41_mask; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_41_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_MPORT_42_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_MPORT_42_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_42_mask; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_42_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_MPORT_43_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_MPORT_43_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_43_mask; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_43_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_MPORT_44_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_MPORT_44_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_44_mask; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_44_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_MPORT_45_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_MPORT_45_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_45_mask; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_45_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_MPORT_46_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_MPORT_46_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_46_mask; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_46_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_MPORT_47_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_MPORT_47_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_47_mask; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_47_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_MPORT_48_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_MPORT_48_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_48_mask; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_48_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_MPORT_49_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_MPORT_49_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_49_mask; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_49_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_MPORT_50_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_MPORT_50_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_50_mask; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_50_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_MPORT_51_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_MPORT_51_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_51_mask; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_51_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_MPORT_52_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_MPORT_52_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_52_mask; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_52_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_MPORT_53_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_MPORT_53_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_53_mask; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_53_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_MPORT_54_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_MPORT_54_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_54_mask; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_54_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_MPORT_55_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_MPORT_55_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_55_mask; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_55_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_MPORT_56_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_MPORT_56_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_56_mask; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_56_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_MPORT_57_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_MPORT_57_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_57_mask; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_57_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_MPORT_58_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_MPORT_58_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_58_mask; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_58_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_MPORT_59_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_MPORT_59_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_59_mask; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_59_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_MPORT_60_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_MPORT_60_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_60_mask; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_60_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_MPORT_61_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_MPORT_61_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_61_mask; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_61_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_MPORT_62_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_MPORT_62_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_62_mask; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_62_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_MPORT_63_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_MPORT_63_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_63_mask; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_63_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_MPORT_64_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_MPORT_64_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_64_mask; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_64_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_MPORT_65_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_MPORT_65_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_65_mask; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_65_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_MPORT_66_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_MPORT_66_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_66_mask; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_66_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_MPORT_67_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_MPORT_67_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_67_mask; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_67_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_MPORT_68_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_MPORT_68_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_68_mask; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_68_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_MPORT_69_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_MPORT_69_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_69_mask; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_69_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_MPORT_70_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_MPORT_70_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_70_mask; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_70_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_MPORT_71_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_MPORT_71_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_71_mask; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_71_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_MPORT_72_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_MPORT_72_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_72_mask; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_72_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_MPORT_73_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_MPORT_73_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_73_mask; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_73_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_MPORT_74_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_MPORT_74_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_74_mask; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_74_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_MPORT_75_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_MPORT_75_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_75_mask; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_75_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_MPORT_76_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_MPORT_76_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_76_mask; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_76_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_MPORT_77_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_MPORT_77_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_77_mask; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_77_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_MPORT_78_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_MPORT_78_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_78_mask; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_78_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_MPORT_79_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_MPORT_79_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_79_mask; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_79_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_MPORT_80_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_MPORT_80_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_80_mask; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_80_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_MPORT_81_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_MPORT_81_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_81_mask; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_81_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_MPORT_82_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_MPORT_82_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_82_mask; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_82_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_MPORT_83_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_MPORT_83_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_83_mask; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_83_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_MPORT_84_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_MPORT_84_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_84_mask; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_84_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_MPORT_85_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_MPORT_85_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_85_mask; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_85_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_MPORT_86_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_MPORT_86_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_86_mask; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_86_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_MPORT_87_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_MPORT_87_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_87_mask; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_87_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_MPORT_88_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_MPORT_88_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_88_mask; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_88_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_MPORT_89_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_MPORT_89_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_89_mask; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_89_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_MPORT_90_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_MPORT_90_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_90_mask; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_90_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_MPORT_91_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_MPORT_91_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_91_mask; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_91_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_MPORT_92_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_MPORT_92_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_92_mask; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_92_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_MPORT_93_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_MPORT_93_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_93_mask; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_93_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_MPORT_94_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_MPORT_94_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_94_mask; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_94_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_MPORT_95_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_MPORT_95_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_95_mask; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_95_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_MPORT_96_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_MPORT_96_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_96_mask; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_96_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_MPORT_97_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_MPORT_97_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_97_mask; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_97_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_MPORT_98_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_MPORT_98_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_98_mask; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_98_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_MPORT_99_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_MPORT_99_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_99_mask; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_99_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_MPORT_100_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_MPORT_100_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_100_mask; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_100_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_MPORT_101_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_MPORT_101_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_101_mask; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_101_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_MPORT_102_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_MPORT_102_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_102_mask; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_102_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_MPORT_103_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_MPORT_103_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_103_mask; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_103_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_MPORT_104_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_MPORT_104_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_104_mask; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_104_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_MPORT_105_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_MPORT_105_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_105_mask; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_105_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_MPORT_106_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_MPORT_106_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_106_mask; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_106_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_MPORT_107_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_MPORT_107_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_107_mask; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_107_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_MPORT_108_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_MPORT_108_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_108_mask; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_108_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_MPORT_109_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_MPORT_109_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_109_mask; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_109_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_MPORT_110_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_MPORT_110_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_110_mask; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_110_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_MPORT_111_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_MPORT_111_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_111_mask; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_111_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_MPORT_112_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_MPORT_112_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_112_mask; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_112_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_MPORT_113_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_MPORT_113_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_113_mask; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_113_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_MPORT_114_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_MPORT_114_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_114_mask; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_114_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_MPORT_115_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_MPORT_115_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_115_mask; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_115_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_MPORT_116_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_MPORT_116_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_116_mask; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_116_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_MPORT_117_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_MPORT_117_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_117_mask; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_117_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_MPORT_118_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_MPORT_118_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_118_mask; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_118_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_MPORT_119_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_MPORT_119_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_119_mask; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_119_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_MPORT_120_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_MPORT_120_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_120_mask; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_120_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_MPORT_121_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_MPORT_121_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_121_mask; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_121_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_MPORT_122_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_MPORT_122_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_122_mask; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_122_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_MPORT_123_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_MPORT_123_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_123_mask; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_123_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_MPORT_124_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_MPORT_124_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_124_mask; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_124_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_MPORT_125_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_MPORT_125_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_125_mask; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_125_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_MPORT_126_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_MPORT_126_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_126_mask; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_126_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_MPORT_127_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_MPORT_127_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_127_mask; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_127_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_MPORT_128_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_MPORT_128_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_128_mask; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_128_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_MPORT_129_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_MPORT_129_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_129_mask; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_129_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_MPORT_130_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_MPORT_130_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_130_mask; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_130_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_MPORT_131_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_MPORT_131_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_131_mask; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_131_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_MPORT_132_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_MPORT_132_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_132_mask; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_132_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_MPORT_133_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_MPORT_133_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_133_mask; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_133_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_MPORT_134_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_MPORT_134_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_134_mask; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_134_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_MPORT_135_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_MPORT_135_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_135_mask; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_135_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_MPORT_136_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_MPORT_136_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_136_mask; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_136_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_MPORT_137_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_MPORT_137_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_137_mask; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_137_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_MPORT_138_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_MPORT_138_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_138_mask; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_138_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_MPORT_139_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_MPORT_139_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_139_mask; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_139_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_MPORT_140_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_MPORT_140_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_140_mask; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_140_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_MPORT_141_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_MPORT_141_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_141_mask; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_141_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_MPORT_142_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_MPORT_142_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_142_mask; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_142_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_MPORT_143_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_MPORT_143_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_143_mask; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_143_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_MPORT_144_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_MPORT_144_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_144_mask; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_144_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_MPORT_145_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_MPORT_145_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_145_mask; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_145_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_MPORT_146_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_MPORT_146_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_146_mask; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_146_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_MPORT_147_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_MPORT_147_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_147_mask; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_147_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_MPORT_148_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_MPORT_148_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_148_mask; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_148_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_MPORT_149_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_MPORT_149_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_149_mask; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_149_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_MPORT_150_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_MPORT_150_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_150_mask; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_150_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_MPORT_151_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_MPORT_151_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_151_mask; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_151_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_MPORT_152_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_MPORT_152_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_152_mask; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_152_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_MPORT_153_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_MPORT_153_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_153_mask; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_153_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_MPORT_154_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_MPORT_154_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_154_mask; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_154_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_MPORT_155_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_MPORT_155_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_155_mask; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_155_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_MPORT_156_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_MPORT_156_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_156_mask; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_156_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_MPORT_157_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_MPORT_157_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_157_mask; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_157_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_MPORT_158_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_MPORT_158_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_158_mask; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_158_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_MPORT_159_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_MPORT_159_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_159_mask; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_159_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_MPORT_160_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_MPORT_160_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_160_mask; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_160_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_MPORT_161_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_MPORT_161_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_161_mask; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_161_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_MPORT_162_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_MPORT_162_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_162_mask; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_162_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_MPORT_163_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_MPORT_163_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_163_mask; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_163_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_MPORT_164_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_MPORT_164_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_164_mask; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_164_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_MPORT_165_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_MPORT_165_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_165_mask; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_165_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_MPORT_166_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_MPORT_166_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_166_mask; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_166_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_MPORT_167_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_MPORT_167_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_167_mask; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_167_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_MPORT_168_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_MPORT_168_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_168_mask; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_168_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_MPORT_169_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_MPORT_169_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_169_mask; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_169_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_MPORT_170_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_MPORT_170_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_170_mask; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_170_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_MPORT_171_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_MPORT_171_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_171_mask; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_171_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_MPORT_172_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_MPORT_172_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_172_mask; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_172_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_MPORT_173_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_MPORT_173_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_173_mask; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_173_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_MPORT_174_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_MPORT_174_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_174_mask; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_174_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_MPORT_175_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_MPORT_175_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_175_mask; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_175_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_MPORT_176_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_MPORT_176_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_176_mask; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_176_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_MPORT_177_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_MPORT_177_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_177_mask; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_177_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_MPORT_178_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_MPORT_178_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_178_mask; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_178_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_MPORT_179_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_MPORT_179_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_179_mask; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_179_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_MPORT_180_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_MPORT_180_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_180_mask; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_180_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_MPORT_181_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_MPORT_181_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_181_mask; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_181_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_MPORT_182_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_MPORT_182_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_182_mask; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_182_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_MPORT_183_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_MPORT_183_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_183_mask; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_183_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_MPORT_184_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_MPORT_184_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_184_mask; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_184_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_MPORT_185_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_MPORT_185_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_185_mask; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_185_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_MPORT_186_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_MPORT_186_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_186_mask; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_186_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_MPORT_187_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_MPORT_187_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_187_mask; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_187_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_MPORT_188_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_MPORT_188_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_188_mask; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_188_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_MPORT_189_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_MPORT_189_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_189_mask; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_189_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_MPORT_190_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_MPORT_190_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_190_mask; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_190_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_MPORT_191_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_MPORT_191_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_191_mask; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_191_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [63:0] rf_MPORT_192_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [7:0] rf_MPORT_192_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_192_mask; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire  rf_MPORT_192_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  wire [1:0] MAX_STEP = io_mixPc ? 2'h3 : 2'h1; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 145:21]
  reg [1:0] set; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 146:20]
  reg [1:0] step; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 147:21]
  reg [1:0] out_set; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 148:24]
  reg [1:0] out_step; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 149:25]
  reg  exec_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 150:24]
  wire  _GEN_0 = io_uart_ctrl_rx_valid | exec_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 151:30 152:13 150:24]
  reg  tx_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 154:22]
  wire  _GEN_1 = io_uart_ctrl_tx_done ? 1'h0 : tx_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 155:29 156:11 154:22]
  reg [255:0] matrix_a_0; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 159:21]
  reg [255:0] matrix_a_1; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 159:21]
  reg [255:0] matrix_a_2; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 159:21]
  reg [255:0] matrix_a_3; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 159:21]
  reg [255:0] matrix_a_4; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 159:21]
  reg [255:0] matrix_a_5; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 159:21]
  reg [255:0] matrix_a_6; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 159:21]
  reg [255:0] matrix_a_7; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 159:21]
  reg [255:0] matrix_b_0; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 160:21]
  reg [255:0] matrix_b_1; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 160:21]
  reg [255:0] matrix_b_2; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 160:21]
  reg [255:0] matrix_b_3; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 160:21]
  reg [255:0] matrix_b_4; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 160:21]
  reg [255:0] matrix_b_5; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 160:21]
  reg [255:0] matrix_b_6; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 160:21]
  reg [255:0] matrix_b_7; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 160:21]
  reg [255:0] matrix_c_0; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 161:21]
  reg [255:0] matrix_c_1; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 161:21]
  reg [255:0] matrix_c_2; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 161:21]
  reg [255:0] matrix_c_3; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 161:21]
  reg [255:0] matrix_c_4; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 161:21]
  reg [255:0] matrix_c_5; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 161:21]
  reg [255:0] matrix_c_6; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 161:21]
  reg [255:0] matrix_c_7; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 161:21]
  wire [1:0] _in_valid_T_2 = set - 2'h1; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 167:58]
  wire  in_valid = out_set == set | out_set == _in_valid_T_2 & out_step > step & exec_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 167:36]
  wire  handshaked = in_valid & io_top_src_ready; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 168:29]
  reg  io_top_src_valid_r; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 169:32]
  reg  io_top_src_bits_ctrl_mixPcMode_r; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 173:46]
  wire  _T_1 = 2'h0 == step; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 212:23]
  wire [63:0] a_tile_v__0 = rf_a_tile_v_0_MPORT_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_a_0_T = {64'h0,a_tile_v__0,128'h0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 216:35]
  wire [63:0] matrix_b_0_tile_v__3 = rf_matrix_b_0_tile_v_3_MPORT_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_0_tile_v__2 = rf_matrix_b_0_tile_v_2_MPORT_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_0_tile_v__1 = rf_matrix_b_0_tile_v_1_MPORT_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_0_tile_v__0 = rf_matrix_b_0_tile_v_0_MPORT_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_b_0_T = {matrix_b_0_tile_v__3,matrix_b_0_tile_v__2,matrix_b_0_tile_v__1,matrix_b_0_tile_v__0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] matrix_c_0_tile_v__3 = rf_matrix_c_0_tile_v_3_MPORT_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_0_tile_v__2 = rf_matrix_c_0_tile_v_2_MPORT_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_0_tile_v__1 = rf_matrix_c_0_tile_v_1_MPORT_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_0_tile_v__0 = rf_matrix_c_0_tile_v_0_MPORT_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_c_0_T = {matrix_c_0_tile_v__3,matrix_c_0_tile_v__2,matrix_c_0_tile_v__1,matrix_c_0_tile_v__0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] a_tile_v_1_2 = rf_a_tile_v_2_MPORT_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] a_tile_v_1_1 = rf_a_tile_v_1_MPORT_1_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] a_tile_v_1_0 = rf_a_tile_v_0_MPORT_1_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] a_1 = {64'h0,a_tile_v_1_2,a_tile_v_1_1,a_tile_v_1_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] matrix_b_0_tile_v_1_3 = rf_matrix_b_0_tile_v_3_MPORT_1_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_0_tile_v_1_2 = rf_matrix_b_0_tile_v_2_MPORT_1_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_0_tile_v_1_1 = rf_matrix_b_0_tile_v_1_MPORT_1_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_0_tile_v_1_0 = rf_matrix_b_0_tile_v_0_MPORT_1_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_b_0_T_1 = {matrix_b_0_tile_v_1_3,matrix_b_0_tile_v_1_2,matrix_b_0_tile_v_1_1,
    matrix_b_0_tile_v_1_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] matrix_c_0_tile_v_1_3 = rf_matrix_c_0_tile_v_3_MPORT_1_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_0_tile_v_1_2 = rf_matrix_c_0_tile_v_2_MPORT_1_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_0_tile_v_1_1 = rf_matrix_c_0_tile_v_1_MPORT_1_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_0_tile_v_1_0 = rf_matrix_c_0_tile_v_0_MPORT_1_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_c_0_T_1 = {matrix_c_0_tile_v_1_3,matrix_c_0_tile_v_1_2,matrix_c_0_tile_v_1_1,
    matrix_c_0_tile_v_1_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire  _GEN_22 = io_mixPc ? 1'h0 : 1'h1; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 214:29 8:15 9:57]
  wire  _T_2 = 2'h1 == step; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 212:23]
  wire [63:0] a_tile_v_2_1 = rf_a_tile_v_1_MPORT_2_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] a_tile_v_2_0 = rf_a_tile_v_0_MPORT_2_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_a_0_T_1 = {a_tile_v_2_1,a_tile_v_2_0,128'h0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 229:35]
  wire [63:0] matrix_b_0_tile_v_2_3 = rf_matrix_b_0_tile_v_3_MPORT_2_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_0_tile_v_2_2 = rf_matrix_b_0_tile_v_2_MPORT_2_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_0_tile_v_2_1 = rf_matrix_b_0_tile_v_1_MPORT_2_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_0_tile_v_2_0 = rf_matrix_b_0_tile_v_0_MPORT_2_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_b_0_T_2 = {matrix_b_0_tile_v_2_3,matrix_b_0_tile_v_2_2,matrix_b_0_tile_v_2_1,
    matrix_b_0_tile_v_2_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] matrix_c_0_tile_v_2_3 = rf_matrix_c_0_tile_v_3_MPORT_2_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_0_tile_v_2_2 = rf_matrix_c_0_tile_v_2_MPORT_2_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_0_tile_v_2_1 = rf_matrix_c_0_tile_v_1_MPORT_2_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_0_tile_v_2_0 = rf_matrix_c_0_tile_v_0_MPORT_2_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_c_0_T_2 = {matrix_c_0_tile_v_2_3,matrix_c_0_tile_v_2_2,matrix_c_0_tile_v_2_1,
    matrix_c_0_tile_v_2_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] a_tile_v_3_2 = rf_a_tile_v_2_MPORT_1_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] a_tile_v_3_1 = rf_a_tile_v_1_MPORT_3_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] a_tile_v_3_0 = rf_a_tile_v_0_MPORT_3_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] a_3 = {64'h0,a_tile_v_3_2,a_tile_v_3_1,a_tile_v_3_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] matrix_b_0_tile_v_3_3 = rf_matrix_b_0_tile_v_3_MPORT_3_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_0_tile_v_3_2 = rf_matrix_b_0_tile_v_2_MPORT_3_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_0_tile_v_3_1 = rf_matrix_b_0_tile_v_1_MPORT_3_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_0_tile_v_3_0 = rf_matrix_b_0_tile_v_0_MPORT_3_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_b_0_T_3 = {matrix_b_0_tile_v_3_3,matrix_b_0_tile_v_3_2,matrix_b_0_tile_v_3_1,
    matrix_b_0_tile_v_3_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] matrix_c_0_tile_v_3_3 = rf_matrix_c_0_tile_v_3_MPORT_3_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_0_tile_v_3_2 = rf_matrix_c_0_tile_v_2_MPORT_3_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_0_tile_v_3_1 = rf_matrix_c_0_tile_v_1_MPORT_3_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_0_tile_v_3_0 = rf_matrix_c_0_tile_v_0_MPORT_3_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_c_0_T_3 = {matrix_c_0_tile_v_3_3,matrix_c_0_tile_v_3_2,matrix_c_0_tile_v_3_1,
    matrix_c_0_tile_v_3_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [255:0] _GEN_36 = io_mixPc ? _matrix_a_0_T_1 : a_3; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 227:30 229:29 234:29]
  wire [255:0] _GEN_37 = io_mixPc ? _matrix_b_0_T_2 : _matrix_b_0_T_3; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 227:30 230:29 235:29]
  wire [255:0] _GEN_42 = io_mixPc ? _matrix_c_0_T_2 : _matrix_c_0_T_3; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 227:30 231:29 236:29]
  wire  _T_3 = 2'h2 == step; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 212:23]
  wire [63:0] a_tile_v_4_0 = rf_a_tile_v_0_MPORT_4_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_a_0_T_2 = {64'h0,a_tile_v_4_0,128'h0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 241:33]
  wire [63:0] matrix_b_0_tile_v_4_3 = rf_matrix_b_0_tile_v_3_MPORT_4_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_0_tile_v_4_2 = rf_matrix_b_0_tile_v_2_MPORT_4_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_0_tile_v_4_1 = rf_matrix_b_0_tile_v_1_MPORT_4_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_0_tile_v_4_0 = rf_matrix_b_0_tile_v_0_MPORT_4_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_b_0_T_4 = {matrix_b_0_tile_v_4_3,matrix_b_0_tile_v_4_2,matrix_b_0_tile_v_4_1,
    matrix_b_0_tile_v_4_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] matrix_c_0_tile_v_4_3 = rf_matrix_c_0_tile_v_3_MPORT_4_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_0_tile_v_4_2 = rf_matrix_c_0_tile_v_2_MPORT_4_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_0_tile_v_4_1 = rf_matrix_c_0_tile_v_1_MPORT_4_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_0_tile_v_4_0 = rf_matrix_c_0_tile_v_0_MPORT_4_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_c_0_T_4 = {matrix_c_0_tile_v_4_3,matrix_c_0_tile_v_4_2,matrix_c_0_tile_v_4_1,
    matrix_c_0_tile_v_4_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire  _T_4 = 2'h3 == step; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 212:23]
  wire [63:0] a_tile_v_5_1 = rf_a_tile_v_1_MPORT_5_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] a_tile_v_5_0 = rf_a_tile_v_0_MPORT_5_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_a_0_T_3 = {a_tile_v_5_1,a_tile_v_5_0,128'h0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 247:33]
  wire [63:0] matrix_b_0_tile_v_5_3 = rf_matrix_b_0_tile_v_3_MPORT_5_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_0_tile_v_5_2 = rf_matrix_b_0_tile_v_2_MPORT_5_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_0_tile_v_5_1 = rf_matrix_b_0_tile_v_1_MPORT_5_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_0_tile_v_5_0 = rf_matrix_b_0_tile_v_0_MPORT_5_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_b_0_T_5 = {matrix_b_0_tile_v_5_3,matrix_b_0_tile_v_5_2,matrix_b_0_tile_v_5_1,
    matrix_b_0_tile_v_5_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] matrix_c_0_tile_v_5_3 = rf_matrix_c_0_tile_v_3_MPORT_5_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_0_tile_v_5_2 = rf_matrix_c_0_tile_v_2_MPORT_5_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_0_tile_v_5_1 = rf_matrix_c_0_tile_v_1_MPORT_5_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_0_tile_v_5_0 = rf_matrix_c_0_tile_v_0_MPORT_5_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_c_0_T_5 = {matrix_c_0_tile_v_5_3,matrix_c_0_tile_v_5_2,matrix_c_0_tile_v_5_1,
    matrix_c_0_tile_v_5_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [255:0] _GEN_51 = 2'h3 == step ? _matrix_a_0_T_3 : matrix_a_0; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 159:21 212:23 247:27]
  wire [255:0] _GEN_56 = 2'h3 == step ? _matrix_b_0_T_5 : matrix_b_0; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 160:21 212:23 248:27]
  wire [255:0] _GEN_61 = 2'h3 == step ? _matrix_c_0_T_5 : matrix_c_0; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 161:21 212:23 249:27]
  wire [255:0] _GEN_66 = 2'h2 == step ? _matrix_a_0_T_2 : _GEN_51; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 212:23 241:27]
  wire [255:0] _GEN_71 = 2'h2 == step ? _matrix_b_0_T_4 : _GEN_56; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 212:23 242:27]
  wire [255:0] _GEN_76 = 2'h2 == step ? _matrix_c_0_T_4 : _GEN_61; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 212:23 243:27]
  wire  _GEN_79 = 2'h2 == step ? 1'h0 : 2'h3 == step; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 212:23 8:15]
  wire  _GEN_120 = 2'h1 == step ? 1'h0 : 2'h2 == step; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 212:23 8:15]
  wire  _GEN_132 = 2'h1 == step ? 1'h0 : _GEN_79; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 212:23 8:15]
  wire  _GEN_144 = 2'h0 == step & io_mixPc; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 212:23 8:15]
  wire  _GEN_159 = 2'h0 == step & _GEN_22; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 212:23 8:15]
  wire  _GEN_173 = 2'h0 == step ? 1'h0 : 2'h1 == step & io_mixPc; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 212:23 8:15]
  wire  _GEN_185 = 2'h0 == step ? 1'h0 : 2'h1 == step & _GEN_22; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 212:23 8:15]
  wire  _GEN_199 = 2'h0 == step ? 1'h0 : _GEN_120; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 212:23 8:15]
  wire  _GEN_211 = 2'h0 == step ? 1'h0 : _GEN_132; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 212:23 8:15]
  wire [63:0] a_tile_v_6_1 = rf_a_tile_v_1_MPORT_6_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] a_tile_v_6_0 = rf_a_tile_v_0_MPORT_6_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_a_0_T_4 = {a_tile_v_6_1,a_tile_v_6_0,128'h0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 258:35]
  wire [63:0] matrix_b_0_tile_v_6_3 = rf_matrix_b_0_tile_v_3_MPORT_6_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_0_tile_v_6_2 = rf_matrix_b_0_tile_v_2_MPORT_6_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_0_tile_v_6_1 = rf_matrix_b_0_tile_v_1_MPORT_6_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_0_tile_v_6_0 = rf_matrix_b_0_tile_v_0_MPORT_6_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_b_0_T_6 = {matrix_b_0_tile_v_6_3,matrix_b_0_tile_v_6_2,matrix_b_0_tile_v_6_1,
    matrix_b_0_tile_v_6_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] matrix_c_0_tile_v_6_3 = rf_matrix_c_0_tile_v_3_MPORT_6_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_0_tile_v_6_2 = rf_matrix_c_0_tile_v_2_MPORT_6_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_0_tile_v_6_1 = rf_matrix_c_0_tile_v_1_MPORT_6_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_0_tile_v_6_0 = rf_matrix_c_0_tile_v_0_MPORT_6_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_c_0_T_6 = {matrix_c_0_tile_v_6_3,matrix_c_0_tile_v_6_2,matrix_c_0_tile_v_6_1,
    matrix_c_0_tile_v_6_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] a_tile_v_7_3 = rf_a_tile_v_3_MPORT_2_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] a_tile_v_7_2 = rf_a_tile_v_2_MPORT_2_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] a_tile_v_7_1 = rf_a_tile_v_1_MPORT_7_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] a_tile_v_7_0 = rf_a_tile_v_0_MPORT_7_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] a_7 = {a_tile_v_7_3,a_tile_v_7_2,a_tile_v_7_1,a_tile_v_7_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] matrix_b_0_tile_v_7_3 = rf_matrix_b_0_tile_v_3_MPORT_7_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_0_tile_v_7_2 = rf_matrix_b_0_tile_v_2_MPORT_7_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_0_tile_v_7_1 = rf_matrix_b_0_tile_v_1_MPORT_7_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_0_tile_v_7_0 = rf_matrix_b_0_tile_v_0_MPORT_7_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_b_0_T_7 = {matrix_b_0_tile_v_7_3,matrix_b_0_tile_v_7_2,matrix_b_0_tile_v_7_1,
    matrix_b_0_tile_v_7_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] matrix_c_0_tile_v_7_3 = rf_matrix_c_0_tile_v_3_MPORT_7_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_0_tile_v_7_2 = rf_matrix_c_0_tile_v_2_MPORT_7_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_0_tile_v_7_1 = rf_matrix_c_0_tile_v_1_MPORT_7_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_0_tile_v_7_0 = rf_matrix_c_0_tile_v_0_MPORT_7_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_c_0_T_7 = {matrix_c_0_tile_v_7_3,matrix_c_0_tile_v_7_2,matrix_c_0_tile_v_7_1,
    matrix_c_0_tile_v_7_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [255:0] _GEN_223 = io_mixPc ? _matrix_a_0_T_4 : a_7; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 256:30 258:29 263:29]
  wire [255:0] _GEN_228 = io_mixPc ? _matrix_b_0_T_6 : _matrix_b_0_T_7; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 256:30 259:29 264:29]
  wire [255:0] _GEN_229 = io_mixPc ? _matrix_c_0_T_6 : _matrix_c_0_T_7; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 256:30 260:29 265:29]
  wire [63:0] a_tile_v_8_1 = rf_a_tile_v_1_MPORT_8_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] a_tile_v_8_0 = rf_a_tile_v_0_MPORT_8_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_a_0_T_5 = {a_tile_v_8_1,a_tile_v_8_0,128'h0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 271:35]
  wire [63:0] matrix_b_0_tile_v_8_3 = rf_matrix_b_0_tile_v_3_MPORT_8_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_0_tile_v_8_2 = rf_matrix_b_0_tile_v_2_MPORT_8_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_0_tile_v_8_1 = rf_matrix_b_0_tile_v_1_MPORT_8_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_0_tile_v_8_0 = rf_matrix_b_0_tile_v_0_MPORT_8_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_b_0_T_8 = {matrix_b_0_tile_v_8_3,matrix_b_0_tile_v_8_2,matrix_b_0_tile_v_8_1,
    matrix_b_0_tile_v_8_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] matrix_c_0_tile_v_8_3 = rf_matrix_c_0_tile_v_3_MPORT_8_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_0_tile_v_8_2 = rf_matrix_c_0_tile_v_2_MPORT_8_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_0_tile_v_8_1 = rf_matrix_c_0_tile_v_1_MPORT_8_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_0_tile_v_8_0 = rf_matrix_c_0_tile_v_0_MPORT_8_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_c_0_T_8 = {matrix_c_0_tile_v_8_3,matrix_c_0_tile_v_8_2,matrix_c_0_tile_v_8_1,
    matrix_c_0_tile_v_8_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] a_tile_v_9_3 = rf_a_tile_v_3_MPORT_3_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] a_tile_v_9_2 = rf_a_tile_v_2_MPORT_3_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] a_tile_v_9_1 = rf_a_tile_v_1_MPORT_9_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] a_tile_v_9_0 = rf_a_tile_v_0_MPORT_9_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] a_9 = {a_tile_v_9_3,a_tile_v_9_2,a_tile_v_9_1,a_tile_v_9_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] matrix_b_0_tile_v_9_3 = rf_matrix_b_0_tile_v_3_MPORT_9_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_0_tile_v_9_2 = rf_matrix_b_0_tile_v_2_MPORT_9_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_0_tile_v_9_1 = rf_matrix_b_0_tile_v_1_MPORT_9_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_0_tile_v_9_0 = rf_matrix_b_0_tile_v_0_MPORT_9_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_b_0_T_9 = {matrix_b_0_tile_v_9_3,matrix_b_0_tile_v_9_2,matrix_b_0_tile_v_9_1,
    matrix_b_0_tile_v_9_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] matrix_c_0_tile_v_9_3 = rf_matrix_c_0_tile_v_3_MPORT_9_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_0_tile_v_9_2 = rf_matrix_c_0_tile_v_2_MPORT_9_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_0_tile_v_9_1 = rf_matrix_c_0_tile_v_1_MPORT_9_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_0_tile_v_9_0 = rf_matrix_c_0_tile_v_0_MPORT_9_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_c_0_T_9 = {matrix_c_0_tile_v_9_3,matrix_c_0_tile_v_9_2,matrix_c_0_tile_v_9_1,
    matrix_c_0_tile_v_9_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [255:0] _GEN_240 = io_mixPc ? _matrix_a_0_T_5 : a_9; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 269:30 271:29 276:29]
  wire [255:0] _GEN_241 = io_mixPc ? _matrix_b_0_T_8 : _matrix_b_0_T_9; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 269:30 272:29 277:29]
  wire [255:0] _GEN_242 = io_mixPc ? _matrix_c_0_T_8 : _matrix_c_0_T_9; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 269:30 273:29 278:29]
  wire [63:0] a_tile_v_10_1 = rf_a_tile_v_1_MPORT_10_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] a_tile_v_10_0 = rf_a_tile_v_0_MPORT_10_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_a_0_T_6 = {a_tile_v_10_1,a_tile_v_10_0,128'h0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 283:33]
  wire [63:0] matrix_b_0_tile_v_10_3 = rf_matrix_b_0_tile_v_3_MPORT_10_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_0_tile_v_10_2 = rf_matrix_b_0_tile_v_2_MPORT_10_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_0_tile_v_10_1 = rf_matrix_b_0_tile_v_1_MPORT_10_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_0_tile_v_10_0 = rf_matrix_b_0_tile_v_0_MPORT_10_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_b_0_T_10 = {matrix_b_0_tile_v_10_3,matrix_b_0_tile_v_10_2,matrix_b_0_tile_v_10_1,
    matrix_b_0_tile_v_10_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] matrix_c_0_tile_v_10_3 = rf_matrix_c_0_tile_v_3_MPORT_10_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_0_tile_v_10_2 = rf_matrix_c_0_tile_v_2_MPORT_10_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_0_tile_v_10_1 = rf_matrix_c_0_tile_v_1_MPORT_10_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_0_tile_v_10_0 = rf_matrix_c_0_tile_v_0_MPORT_10_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_c_0_T_10 = {matrix_c_0_tile_v_10_3,matrix_c_0_tile_v_10_2,matrix_c_0_tile_v_10_1,
    matrix_c_0_tile_v_10_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] a_tile_v_11_1 = rf_a_tile_v_1_MPORT_11_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] a_tile_v_11_0 = rf_a_tile_v_0_MPORT_11_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_a_0_T_7 = {a_tile_v_11_1,a_tile_v_11_0,128'h0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 289:33]
  wire [63:0] matrix_b_0_tile_v_11_3 = rf_matrix_b_0_tile_v_3_MPORT_11_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_0_tile_v_11_2 = rf_matrix_b_0_tile_v_2_MPORT_11_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_0_tile_v_11_1 = rf_matrix_b_0_tile_v_1_MPORT_11_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_0_tile_v_11_0 = rf_matrix_b_0_tile_v_0_MPORT_11_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_b_0_T_11 = {matrix_b_0_tile_v_11_3,matrix_b_0_tile_v_11_2,matrix_b_0_tile_v_11_1,
    matrix_b_0_tile_v_11_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] matrix_c_0_tile_v_11_3 = rf_matrix_c_0_tile_v_3_MPORT_11_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_0_tile_v_11_2 = rf_matrix_c_0_tile_v_2_MPORT_11_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_0_tile_v_11_1 = rf_matrix_c_0_tile_v_1_MPORT_11_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_0_tile_v_11_0 = rf_matrix_c_0_tile_v_0_MPORT_11_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_c_0_T_11 = {matrix_c_0_tile_v_11_3,matrix_c_0_tile_v_11_2,matrix_c_0_tile_v_11_1,
    matrix_c_0_tile_v_11_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [255:0] _GEN_247 = _T_4 ? _matrix_a_0_T_7 : matrix_a_0; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 159:21 254:24 289:27]
  wire [255:0] _GEN_252 = _T_4 ? _matrix_b_0_T_11 : matrix_b_0; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 160:21 254:24 290:27]
  wire [255:0] _GEN_257 = _T_4 ? _matrix_c_0_T_11 : matrix_c_0; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 161:21 254:24 291:27]
  wire [255:0] _GEN_262 = _T_3 ? _matrix_a_0_T_6 : _GEN_247; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 254:24 283:27]
  wire [255:0] _GEN_267 = _T_3 ? _matrix_b_0_T_10 : _GEN_252; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 254:24 284:27]
  wire [255:0] _GEN_272 = _T_3 ? _matrix_c_0_T_10 : _GEN_257; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 254:24 285:27]
  wire [255:0] _GEN_289 = _T_2 ? _GEN_240 : _GEN_262; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 254:24]
  wire [255:0] _GEN_294 = _T_2 ? _GEN_241 : _GEN_267; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 254:24]
  wire [255:0] _GEN_299 = _T_2 ? _GEN_242 : _GEN_272; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 254:24]
  wire [63:0] a_tile_v_12_1 = rf_a_tile_v_1_MPORT_12_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] a_tile_v_12_0 = rf_a_tile_v_0_MPORT_12_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_a_0_T_8 = {a_tile_v_12_1,a_tile_v_12_0,128'h0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 300:35]
  wire [63:0] matrix_b_0_tile_v_12_3 = rf_matrix_b_0_tile_v_3_MPORT_12_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_0_tile_v_12_2 = rf_matrix_b_0_tile_v_2_MPORT_12_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_0_tile_v_12_1 = rf_matrix_b_0_tile_v_1_MPORT_12_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_0_tile_v_12_0 = rf_matrix_b_0_tile_v_0_MPORT_12_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_b_0_T_12 = {matrix_b_0_tile_v_12_3,matrix_b_0_tile_v_12_2,matrix_b_0_tile_v_12_1,
    matrix_b_0_tile_v_12_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] matrix_c_0_tile_v_12_3 = rf_matrix_c_0_tile_v_3_MPORT_12_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_0_tile_v_12_2 = rf_matrix_c_0_tile_v_2_MPORT_12_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_0_tile_v_12_1 = rf_matrix_c_0_tile_v_1_MPORT_12_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_0_tile_v_12_0 = rf_matrix_c_0_tile_v_0_MPORT_12_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_c_0_T_12 = {matrix_c_0_tile_v_12_3,matrix_c_0_tile_v_12_2,matrix_c_0_tile_v_12_1,
    matrix_c_0_tile_v_12_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] a_tile_v_13_3 = rf_a_tile_v_3_MPORT_4_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] a_tile_v_13_2 = rf_a_tile_v_2_MPORT_4_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] a_tile_v_13_1 = rf_a_tile_v_1_MPORT_13_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] a_tile_v_13_0 = rf_a_tile_v_0_MPORT_13_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] a_13 = {a_tile_v_13_3,a_tile_v_13_2,a_tile_v_13_1,a_tile_v_13_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] matrix_b_0_tile_v_13_3 = rf_matrix_b_0_tile_v_3_MPORT_13_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_0_tile_v_13_2 = rf_matrix_b_0_tile_v_2_MPORT_13_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_0_tile_v_13_1 = rf_matrix_b_0_tile_v_1_MPORT_13_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_0_tile_v_13_0 = rf_matrix_b_0_tile_v_0_MPORT_13_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_b_0_T_13 = {matrix_b_0_tile_v_13_3,matrix_b_0_tile_v_13_2,matrix_b_0_tile_v_13_1,
    matrix_b_0_tile_v_13_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] matrix_c_0_tile_v_13_3 = rf_matrix_c_0_tile_v_3_MPORT_13_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_0_tile_v_13_2 = rf_matrix_c_0_tile_v_2_MPORT_13_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_0_tile_v_13_1 = rf_matrix_c_0_tile_v_1_MPORT_13_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_0_tile_v_13_0 = rf_matrix_c_0_tile_v_0_MPORT_13_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_c_0_T_13 = {matrix_c_0_tile_v_13_3,matrix_c_0_tile_v_13_2,matrix_c_0_tile_v_13_1,
    matrix_c_0_tile_v_13_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [255:0] _GEN_419 = io_mixPc ? _matrix_a_0_T_8 : a_13; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 298:30 300:29 305:29]
  wire [255:0] _GEN_424 = io_mixPc ? _matrix_b_0_T_12 : _matrix_b_0_T_13; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 298:30 301:29 306:29]
  wire [255:0] _GEN_425 = io_mixPc ? _matrix_c_0_T_12 : _matrix_c_0_T_13; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 298:30 302:29 307:29]
  wire [63:0] a_tile_v_14_1 = rf_a_tile_v_1_MPORT_14_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] a_tile_v_14_0 = rf_a_tile_v_0_MPORT_14_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_a_0_T_9 = {a_tile_v_14_1,a_tile_v_14_0,128'h0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 313:35]
  wire [63:0] matrix_b_0_tile_v_14_3 = rf_matrix_b_0_tile_v_3_MPORT_14_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_0_tile_v_14_2 = rf_matrix_b_0_tile_v_2_MPORT_14_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_0_tile_v_14_1 = rf_matrix_b_0_tile_v_1_MPORT_14_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_0_tile_v_14_0 = rf_matrix_b_0_tile_v_0_MPORT_14_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_b_0_T_14 = {matrix_b_0_tile_v_14_3,matrix_b_0_tile_v_14_2,matrix_b_0_tile_v_14_1,
    matrix_b_0_tile_v_14_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] matrix_c_0_tile_v_14_3 = rf_matrix_c_0_tile_v_3_MPORT_14_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_0_tile_v_14_2 = rf_matrix_c_0_tile_v_2_MPORT_14_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_0_tile_v_14_1 = rf_matrix_c_0_tile_v_1_MPORT_14_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_0_tile_v_14_0 = rf_matrix_c_0_tile_v_0_MPORT_14_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_c_0_T_14 = {matrix_c_0_tile_v_14_3,matrix_c_0_tile_v_14_2,matrix_c_0_tile_v_14_1,
    matrix_c_0_tile_v_14_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] a_tile_v_15_3 = rf_a_tile_v_3_MPORT_5_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] a_tile_v_15_2 = rf_a_tile_v_2_MPORT_5_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] a_tile_v_15_1 = rf_a_tile_v_1_MPORT_15_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] a_tile_v_15_0 = rf_a_tile_v_0_MPORT_15_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] a_15 = {a_tile_v_15_3,a_tile_v_15_2,a_tile_v_15_1,a_tile_v_15_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] matrix_b_0_tile_v_15_3 = rf_matrix_b_0_tile_v_3_MPORT_15_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_0_tile_v_15_2 = rf_matrix_b_0_tile_v_2_MPORT_15_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_0_tile_v_15_1 = rf_matrix_b_0_tile_v_1_MPORT_15_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_0_tile_v_15_0 = rf_matrix_b_0_tile_v_0_MPORT_15_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_b_0_T_15 = {matrix_b_0_tile_v_15_3,matrix_b_0_tile_v_15_2,matrix_b_0_tile_v_15_1,
    matrix_b_0_tile_v_15_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] matrix_c_0_tile_v_15_3 = rf_matrix_c_0_tile_v_3_MPORT_15_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_0_tile_v_15_2 = rf_matrix_c_0_tile_v_2_MPORT_15_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_0_tile_v_15_1 = rf_matrix_c_0_tile_v_1_MPORT_15_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_0_tile_v_15_0 = rf_matrix_c_0_tile_v_0_MPORT_15_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_c_0_T_15 = {matrix_c_0_tile_v_15_3,matrix_c_0_tile_v_15_2,matrix_c_0_tile_v_15_1,
    matrix_c_0_tile_v_15_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [255:0] _GEN_436 = io_mixPc ? _matrix_a_0_T_9 : a_15; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 311:30 313:29 318:29]
  wire [255:0] _GEN_437 = io_mixPc ? _matrix_b_0_T_14 : _matrix_b_0_T_15; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 311:30 314:29 319:29]
  wire [255:0] _GEN_438 = io_mixPc ? _matrix_c_0_T_14 : _matrix_c_0_T_15; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 311:30 315:29 320:29]
  wire [63:0] a_tile_v_16_1 = rf_a_tile_v_1_MPORT_16_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] a_tile_v_16_0 = rf_a_tile_v_0_MPORT_16_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_a_0_T_10 = {a_tile_v_16_1,a_tile_v_16_0,128'h0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 325:33]
  wire [63:0] matrix_b_0_tile_v_16_3 = rf_matrix_b_0_tile_v_3_MPORT_16_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_0_tile_v_16_2 = rf_matrix_b_0_tile_v_2_MPORT_16_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_0_tile_v_16_1 = rf_matrix_b_0_tile_v_1_MPORT_16_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_0_tile_v_16_0 = rf_matrix_b_0_tile_v_0_MPORT_16_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_b_0_T_16 = {matrix_b_0_tile_v_16_3,matrix_b_0_tile_v_16_2,matrix_b_0_tile_v_16_1,
    matrix_b_0_tile_v_16_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] matrix_c_0_tile_v_16_3 = rf_matrix_c_0_tile_v_3_MPORT_16_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_0_tile_v_16_2 = rf_matrix_c_0_tile_v_2_MPORT_16_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_0_tile_v_16_1 = rf_matrix_c_0_tile_v_1_MPORT_16_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_0_tile_v_16_0 = rf_matrix_c_0_tile_v_0_MPORT_16_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_c_0_T_16 = {matrix_c_0_tile_v_16_3,matrix_c_0_tile_v_16_2,matrix_c_0_tile_v_16_1,
    matrix_c_0_tile_v_16_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] a_tile_v_17_1 = rf_a_tile_v_1_MPORT_17_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] a_tile_v_17_0 = rf_a_tile_v_0_MPORT_17_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_a_0_T_11 = {a_tile_v_17_1,a_tile_v_17_0,128'h0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 331:33]
  wire [63:0] matrix_b_0_tile_v_17_3 = rf_matrix_b_0_tile_v_3_MPORT_17_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_0_tile_v_17_2 = rf_matrix_b_0_tile_v_2_MPORT_17_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_0_tile_v_17_1 = rf_matrix_b_0_tile_v_1_MPORT_17_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_0_tile_v_17_0 = rf_matrix_b_0_tile_v_0_MPORT_17_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_b_0_T_17 = {matrix_b_0_tile_v_17_3,matrix_b_0_tile_v_17_2,matrix_b_0_tile_v_17_1,
    matrix_b_0_tile_v_17_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] matrix_c_0_tile_v_17_3 = rf_matrix_c_0_tile_v_3_MPORT_17_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_0_tile_v_17_2 = rf_matrix_c_0_tile_v_2_MPORT_17_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_0_tile_v_17_1 = rf_matrix_c_0_tile_v_1_MPORT_17_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_0_tile_v_17_0 = rf_matrix_c_0_tile_v_0_MPORT_17_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_c_0_T_17 = {matrix_c_0_tile_v_17_3,matrix_c_0_tile_v_17_2,matrix_c_0_tile_v_17_1,
    matrix_c_0_tile_v_17_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [255:0] _GEN_443 = _T_4 ? _matrix_a_0_T_11 : matrix_a_0; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 159:21 296:24 331:27]
  wire [255:0] _GEN_448 = _T_4 ? _matrix_b_0_T_17 : matrix_b_0; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 160:21 296:24 332:27]
  wire [255:0] _GEN_453 = _T_4 ? _matrix_c_0_T_17 : matrix_c_0; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 161:21 296:24 333:27]
  wire [255:0] _GEN_458 = _T_3 ? _matrix_a_0_T_10 : _GEN_443; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 296:24 325:27]
  wire [255:0] _GEN_463 = _T_3 ? _matrix_b_0_T_16 : _GEN_448; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 296:24 326:27]
  wire [255:0] _GEN_468 = _T_3 ? _matrix_c_0_T_16 : _GEN_453; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 296:24 327:27]
  wire [255:0] _GEN_485 = _T_2 ? _GEN_436 : _GEN_458; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 296:24]
  wire [255:0] _GEN_490 = _T_2 ? _GEN_437 : _GEN_463; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 296:24]
  wire [255:0] _GEN_495 = _T_2 ? _GEN_438 : _GEN_468; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 296:24]
  wire [255:0] _GEN_538 = _T_1 ? _GEN_419 : _GEN_485; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 296:24]
  wire [255:0] _GEN_543 = _T_1 ? _GEN_424 : _GEN_490; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 296:24]
  wire [255:0] _GEN_548 = _T_1 ? _GEN_425 : _GEN_495; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 296:24]
  wire [63:0] a_tile_v_18_1 = rf_a_tile_v_1_MPORT_18_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] a_tile_v_18_0 = rf_a_tile_v_0_MPORT_18_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_a_0_T_12 = {a_tile_v_18_1,a_tile_v_18_0,128'h0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 342:35]
  wire [63:0] matrix_b_0_tile_v_18_3 = rf_matrix_b_0_tile_v_3_MPORT_18_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_0_tile_v_18_2 = rf_matrix_b_0_tile_v_2_MPORT_18_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_0_tile_v_18_1 = rf_matrix_b_0_tile_v_1_MPORT_18_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_0_tile_v_18_0 = rf_matrix_b_0_tile_v_0_MPORT_18_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_b_0_T_18 = {matrix_b_0_tile_v_18_3,matrix_b_0_tile_v_18_2,matrix_b_0_tile_v_18_1,
    matrix_b_0_tile_v_18_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] matrix_c_0_tile_v_18_3 = rf_matrix_c_0_tile_v_3_MPORT_18_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_0_tile_v_18_2 = rf_matrix_c_0_tile_v_2_MPORT_18_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_0_tile_v_18_1 = rf_matrix_c_0_tile_v_1_MPORT_18_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_0_tile_v_18_0 = rf_matrix_c_0_tile_v_0_MPORT_18_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_c_0_T_18 = {matrix_c_0_tile_v_18_3,matrix_c_0_tile_v_18_2,matrix_c_0_tile_v_18_1,
    matrix_c_0_tile_v_18_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] a_tile_v_19_3 = rf_a_tile_v_3_MPORT_6_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] a_tile_v_19_2 = rf_a_tile_v_2_MPORT_6_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] a_tile_v_19_1 = rf_a_tile_v_1_MPORT_19_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] a_tile_v_19_0 = rf_a_tile_v_0_MPORT_19_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] a_19 = {a_tile_v_19_3,a_tile_v_19_2,a_tile_v_19_1,a_tile_v_19_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] matrix_b_0_tile_v_19_3 = rf_matrix_b_0_tile_v_3_MPORT_19_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_0_tile_v_19_2 = rf_matrix_b_0_tile_v_2_MPORT_19_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_0_tile_v_19_1 = rf_matrix_b_0_tile_v_1_MPORT_19_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_0_tile_v_19_0 = rf_matrix_b_0_tile_v_0_MPORT_19_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_b_0_T_19 = {matrix_b_0_tile_v_19_3,matrix_b_0_tile_v_19_2,matrix_b_0_tile_v_19_1,
    matrix_b_0_tile_v_19_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] matrix_c_0_tile_v_19_3 = rf_matrix_c_0_tile_v_3_MPORT_19_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_0_tile_v_19_2 = rf_matrix_c_0_tile_v_2_MPORT_19_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_0_tile_v_19_1 = rf_matrix_c_0_tile_v_1_MPORT_19_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_0_tile_v_19_0 = rf_matrix_c_0_tile_v_0_MPORT_19_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_c_0_T_19 = {matrix_c_0_tile_v_19_3,matrix_c_0_tile_v_19_2,matrix_c_0_tile_v_19_1,
    matrix_c_0_tile_v_19_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [255:0] _GEN_615 = io_mixPc ? _matrix_a_0_T_12 : a_19; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 340:30 342:29 347:29]
  wire [255:0] _GEN_620 = io_mixPc ? _matrix_b_0_T_18 : _matrix_b_0_T_19; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 340:30 343:29 348:29]
  wire [255:0] _GEN_621 = io_mixPc ? _matrix_c_0_T_18 : _matrix_c_0_T_19; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 340:30 344:29 349:29]
  wire [63:0] a_tile_v_20_1 = rf_a_tile_v_1_MPORT_20_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] a_tile_v_20_0 = rf_a_tile_v_0_MPORT_20_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_a_0_T_13 = {a_tile_v_20_1,a_tile_v_20_0,128'h0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 355:35]
  wire [63:0] matrix_b_0_tile_v_20_3 = rf_matrix_b_0_tile_v_3_MPORT_20_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_0_tile_v_20_2 = rf_matrix_b_0_tile_v_2_MPORT_20_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_0_tile_v_20_1 = rf_matrix_b_0_tile_v_1_MPORT_20_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_0_tile_v_20_0 = rf_matrix_b_0_tile_v_0_MPORT_20_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_b_0_T_20 = {matrix_b_0_tile_v_20_3,matrix_b_0_tile_v_20_2,matrix_b_0_tile_v_20_1,
    matrix_b_0_tile_v_20_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] matrix_c_0_tile_v_20_3 = rf_matrix_c_0_tile_v_3_MPORT_20_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_0_tile_v_20_2 = rf_matrix_c_0_tile_v_2_MPORT_20_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_0_tile_v_20_1 = rf_matrix_c_0_tile_v_1_MPORT_20_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_0_tile_v_20_0 = rf_matrix_c_0_tile_v_0_MPORT_20_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_c_0_T_20 = {matrix_c_0_tile_v_20_3,matrix_c_0_tile_v_20_2,matrix_c_0_tile_v_20_1,
    matrix_c_0_tile_v_20_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] a_tile_v_21_3 = rf_a_tile_v_3_MPORT_7_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] a_tile_v_21_2 = rf_a_tile_v_2_MPORT_7_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] a_tile_v_21_1 = rf_a_tile_v_1_MPORT_21_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] a_tile_v_21_0 = rf_a_tile_v_0_MPORT_21_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] a_21 = {a_tile_v_21_3,a_tile_v_21_2,a_tile_v_21_1,a_tile_v_21_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] matrix_b_0_tile_v_21_3 = rf_matrix_b_0_tile_v_3_MPORT_21_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_0_tile_v_21_2 = rf_matrix_b_0_tile_v_2_MPORT_21_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_0_tile_v_21_1 = rf_matrix_b_0_tile_v_1_MPORT_21_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_0_tile_v_21_0 = rf_matrix_b_0_tile_v_0_MPORT_21_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_b_0_T_21 = {matrix_b_0_tile_v_21_3,matrix_b_0_tile_v_21_2,matrix_b_0_tile_v_21_1,
    matrix_b_0_tile_v_21_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] matrix_c_0_tile_v_21_3 = rf_matrix_c_0_tile_v_3_MPORT_21_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_0_tile_v_21_2 = rf_matrix_c_0_tile_v_2_MPORT_21_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_0_tile_v_21_1 = rf_matrix_c_0_tile_v_1_MPORT_21_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_0_tile_v_21_0 = rf_matrix_c_0_tile_v_0_MPORT_21_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_c_0_T_21 = {matrix_c_0_tile_v_21_3,matrix_c_0_tile_v_21_2,matrix_c_0_tile_v_21_1,
    matrix_c_0_tile_v_21_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [255:0] _GEN_632 = io_mixPc ? _matrix_a_0_T_13 : a_21; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 353:30 355:29 360:29]
  wire [255:0] _GEN_633 = io_mixPc ? _matrix_b_0_T_20 : _matrix_b_0_T_21; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 353:30 356:29 361:29]
  wire [255:0] _GEN_634 = io_mixPc ? _matrix_c_0_T_20 : _matrix_c_0_T_21; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 353:30 357:29 362:29]
  wire [63:0] a_tile_v_22_1 = rf_a_tile_v_1_MPORT_22_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] a_tile_v_22_0 = rf_a_tile_v_0_MPORT_22_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_a_0_T_14 = {a_tile_v_22_1,a_tile_v_22_0,128'h0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 367:33]
  wire [63:0] matrix_b_0_tile_v_22_3 = rf_matrix_b_0_tile_v_3_MPORT_22_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_0_tile_v_22_2 = rf_matrix_b_0_tile_v_2_MPORT_22_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_0_tile_v_22_1 = rf_matrix_b_0_tile_v_1_MPORT_22_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_0_tile_v_22_0 = rf_matrix_b_0_tile_v_0_MPORT_22_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_b_0_T_22 = {matrix_b_0_tile_v_22_3,matrix_b_0_tile_v_22_2,matrix_b_0_tile_v_22_1,
    matrix_b_0_tile_v_22_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] matrix_c_0_tile_v_22_3 = rf_matrix_c_0_tile_v_3_MPORT_22_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_0_tile_v_22_2 = rf_matrix_c_0_tile_v_2_MPORT_22_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_0_tile_v_22_1 = rf_matrix_c_0_tile_v_1_MPORT_22_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_0_tile_v_22_0 = rf_matrix_c_0_tile_v_0_MPORT_22_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_c_0_T_22 = {matrix_c_0_tile_v_22_3,matrix_c_0_tile_v_22_2,matrix_c_0_tile_v_22_1,
    matrix_c_0_tile_v_22_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] a_tile_v_23_1 = rf_a_tile_v_1_MPORT_23_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] a_tile_v_23_0 = rf_a_tile_v_0_MPORT_23_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_a_0_T_15 = {a_tile_v_23_1,a_tile_v_23_0,128'h0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 373:33]
  wire [63:0] matrix_b_0_tile_v_23_3 = rf_matrix_b_0_tile_v_3_MPORT_23_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_0_tile_v_23_2 = rf_matrix_b_0_tile_v_2_MPORT_23_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_0_tile_v_23_1 = rf_matrix_b_0_tile_v_1_MPORT_23_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_0_tile_v_23_0 = rf_matrix_b_0_tile_v_0_MPORT_23_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_b_0_T_23 = {matrix_b_0_tile_v_23_3,matrix_b_0_tile_v_23_2,matrix_b_0_tile_v_23_1,
    matrix_b_0_tile_v_23_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] matrix_c_0_tile_v_23_3 = rf_matrix_c_0_tile_v_3_MPORT_23_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_0_tile_v_23_2 = rf_matrix_c_0_tile_v_2_MPORT_23_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_0_tile_v_23_1 = rf_matrix_c_0_tile_v_1_MPORT_23_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_0_tile_v_23_0 = rf_matrix_c_0_tile_v_0_MPORT_23_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_c_0_T_23 = {matrix_c_0_tile_v_23_3,matrix_c_0_tile_v_23_2,matrix_c_0_tile_v_23_1,
    matrix_c_0_tile_v_23_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [255:0] _GEN_639 = _T_4 ? _matrix_a_0_T_15 : matrix_a_0; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 159:21 338:24 373:27]
  wire [255:0] _GEN_644 = _T_4 ? _matrix_b_0_T_23 : matrix_b_0; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 160:21 338:24 374:27]
  wire [255:0] _GEN_649 = _T_4 ? _matrix_c_0_T_23 : matrix_c_0; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 161:21 338:24 375:27]
  wire [255:0] _GEN_654 = _T_3 ? _matrix_a_0_T_14 : _GEN_639; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 338:24 367:27]
  wire [255:0] _GEN_659 = _T_3 ? _matrix_b_0_T_22 : _GEN_644; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 338:24 368:27]
  wire [255:0] _GEN_664 = _T_3 ? _matrix_c_0_T_22 : _GEN_649; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 338:24 369:27]
  wire [255:0] _GEN_681 = _T_2 ? _GEN_632 : _GEN_654; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 338:24]
  wire [255:0] _GEN_686 = _T_2 ? _GEN_633 : _GEN_659; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 338:24]
  wire [255:0] _GEN_691 = _T_2 ? _GEN_634 : _GEN_664; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 338:24]
  wire [255:0] _GEN_734 = _T_1 ? _GEN_615 : _GEN_681; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 338:24]
  wire [255:0] _GEN_739 = _T_1 ? _GEN_620 : _GEN_686; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 338:24]
  wire [255:0] _GEN_744 = _T_1 ? _GEN_621 : _GEN_691; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 338:24]
  wire [255:0] _GEN_813 = 2'h3 == set ? _GEN_734 : matrix_a_0; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 210:18 159:21]
  wire [255:0] _GEN_818 = 2'h3 == set ? _GEN_739 : matrix_b_0; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 210:18 160:21]
  wire [255:0] _GEN_823 = 2'h3 == set ? _GEN_744 : matrix_c_0; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 210:18 161:21]
  wire  _GEN_969 = 2'h2 == set ? 1'h0 : 2'h3 == set & _GEN_144; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 210:18 8:15]
  wire  _GEN_981 = 2'h2 == set ? 1'h0 : 2'h3 == set & _GEN_159; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 210:18 8:15]
  wire  _GEN_995 = 2'h2 == set ? 1'h0 : 2'h3 == set & _GEN_173; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 210:18 8:15]
  wire  _GEN_1007 = 2'h2 == set ? 1'h0 : 2'h3 == set & _GEN_185; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 210:18 8:15]
  wire  _GEN_1021 = 2'h2 == set ? 1'h0 : 2'h3 == set & _GEN_199; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 210:18 8:15]
  wire  _GEN_1033 = 2'h2 == set ? 1'h0 : 2'h3 == set & _GEN_211; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 210:18 8:15]
  wire  _GEN_1124 = 2'h1 == set ? 1'h0 : 2'h2 == set & _GEN_144; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 210:18 8:15]
  wire  _GEN_1136 = 2'h1 == set ? 1'h0 : 2'h2 == set & _GEN_159; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 210:18 8:15]
  wire  _GEN_1150 = 2'h1 == set ? 1'h0 : 2'h2 == set & _GEN_173; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 210:18 8:15]
  wire  _GEN_1162 = 2'h1 == set ? 1'h0 : 2'h2 == set & _GEN_185; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 210:18 8:15]
  wire  _GEN_1176 = 2'h1 == set ? 1'h0 : 2'h2 == set & _GEN_199; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 210:18 8:15]
  wire  _GEN_1188 = 2'h1 == set ? 1'h0 : 2'h2 == set & _GEN_211; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 210:18 8:15]
  wire  _GEN_1200 = 2'h1 == set ? 1'h0 : _GEN_969; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 210:18 8:15]
  wire  _GEN_1212 = 2'h1 == set ? 1'h0 : _GEN_981; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 210:18 8:15]
  wire  _GEN_1226 = 2'h1 == set ? 1'h0 : _GEN_995; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 210:18 8:15]
  wire  _GEN_1238 = 2'h1 == set ? 1'h0 : _GEN_1007; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 210:18 8:15]
  wire  _GEN_1252 = 2'h1 == set ? 1'h0 : _GEN_1021; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 210:18 8:15]
  wire  _GEN_1264 = 2'h1 == set ? 1'h0 : _GEN_1033; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 210:18 8:15]
  wire  _GEN_1276 = 2'h0 == set & _GEN_144; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 210:18 8:15]
  wire  _GEN_1291 = 2'h0 == set & _GEN_159; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 210:18 8:15]
  wire  _GEN_1305 = 2'h0 == set & _GEN_173; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 210:18 8:15]
  wire  _GEN_1317 = 2'h0 == set & _GEN_185; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 210:18 8:15]
  wire  _GEN_1331 = 2'h0 == set & _GEN_199; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 210:18 8:15]
  wire  _GEN_1343 = 2'h0 == set & _GEN_211; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 210:18 8:15]
  wire  _GEN_1355 = 2'h0 == set ? 1'h0 : 2'h1 == set & _GEN_144; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 210:18 8:15]
  wire  _GEN_1367 = 2'h0 == set ? 1'h0 : 2'h1 == set & _GEN_159; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 210:18 8:15]
  wire  _GEN_1381 = 2'h0 == set ? 1'h0 : 2'h1 == set & _GEN_173; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 210:18 8:15]
  wire  _GEN_1393 = 2'h0 == set ? 1'h0 : 2'h1 == set & _GEN_185; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 210:18 8:15]
  wire  _GEN_1407 = 2'h0 == set ? 1'h0 : 2'h1 == set & _GEN_199; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 210:18 8:15]
  wire  _GEN_1419 = 2'h0 == set ? 1'h0 : 2'h1 == set & _GEN_211; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 210:18 8:15]
  wire  _GEN_1431 = 2'h0 == set ? 1'h0 : _GEN_1124; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 210:18 8:15]
  wire  _GEN_1443 = 2'h0 == set ? 1'h0 : _GEN_1136; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 210:18 8:15]
  wire  _GEN_1457 = 2'h0 == set ? 1'h0 : _GEN_1150; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 210:18 8:15]
  wire  _GEN_1469 = 2'h0 == set ? 1'h0 : _GEN_1162; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 210:18 8:15]
  wire  _GEN_1483 = 2'h0 == set ? 1'h0 : _GEN_1176; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 210:18 8:15]
  wire  _GEN_1495 = 2'h0 == set ? 1'h0 : _GEN_1188; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 210:18 8:15]
  wire  _GEN_1507 = 2'h0 == set ? 1'h0 : _GEN_1200; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 210:18 8:15]
  wire  _GEN_1519 = 2'h0 == set ? 1'h0 : _GEN_1212; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 210:18 8:15]
  wire  _GEN_1533 = 2'h0 == set ? 1'h0 : _GEN_1226; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 210:18 8:15]
  wire  _GEN_1545 = 2'h0 == set ? 1'h0 : _GEN_1238; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 210:18 8:15]
  wire  _GEN_1559 = 2'h0 == set ? 1'h0 : _GEN_1252; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 210:18 8:15]
  wire  _GEN_1571 = 2'h0 == set ? 1'h0 : _GEN_1264; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 210:18 8:15]
  wire [63:0] a_tile_v_24_1 = rf_a_tile_v_1_MPORT_24_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] a_tile_v_24_0 = rf_a_tile_v_0_MPORT_24_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_a_1_T = {a_tile_v_24_1,a_tile_v_24_0,128'h0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 216:35]
  wire [63:0] matrix_b_1_tile_v__3 = rf_matrix_b_1_tile_v_3_MPORT_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_1_tile_v__2 = rf_matrix_b_1_tile_v_2_MPORT_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_1_tile_v__1 = rf_matrix_b_1_tile_v_1_MPORT_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_1_tile_v__0 = rf_matrix_b_1_tile_v_0_MPORT_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_b_1_T = {matrix_b_1_tile_v__3,matrix_b_1_tile_v__2,matrix_b_1_tile_v__1,matrix_b_1_tile_v__0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] matrix_c_1_tile_v__3 = rf_matrix_c_1_tile_v_3_MPORT_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_1_tile_v__2 = rf_matrix_c_1_tile_v_2_MPORT_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_1_tile_v__1 = rf_matrix_c_1_tile_v_1_MPORT_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_1_tile_v__0 = rf_matrix_c_1_tile_v_0_MPORT_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_c_1_T = {matrix_c_1_tile_v__3,matrix_c_1_tile_v__2,matrix_c_1_tile_v__1,matrix_c_1_tile_v__0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] a_tile_v_25_3 = rf_a_tile_v_3_MPORT_8_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] a_tile_v_25_2 = rf_a_tile_v_2_MPORT_8_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] a_tile_v_25_1 = rf_a_tile_v_1_MPORT_25_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] a_tile_v_25_0 = rf_a_tile_v_0_MPORT_25_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] a_25 = {a_tile_v_25_3,a_tile_v_25_2,a_tile_v_25_1,a_tile_v_25_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] matrix_b_1_tile_v_1_3 = rf_matrix_b_1_tile_v_3_MPORT_1_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_1_tile_v_1_2 = rf_matrix_b_1_tile_v_2_MPORT_1_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_1_tile_v_1_1 = rf_matrix_b_1_tile_v_1_MPORT_1_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_1_tile_v_1_0 = rf_matrix_b_1_tile_v_0_MPORT_1_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_b_1_T_1 = {matrix_b_1_tile_v_1_3,matrix_b_1_tile_v_1_2,matrix_b_1_tile_v_1_1,
    matrix_b_1_tile_v_1_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] matrix_c_1_tile_v_1_3 = rf_matrix_c_1_tile_v_3_MPORT_1_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_1_tile_v_1_2 = rf_matrix_c_1_tile_v_2_MPORT_1_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_1_tile_v_1_1 = rf_matrix_c_1_tile_v_1_MPORT_1_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_1_tile_v_1_0 = rf_matrix_c_1_tile_v_0_MPORT_1_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_c_1_T_1 = {matrix_c_1_tile_v_1_3,matrix_c_1_tile_v_1_2,matrix_c_1_tile_v_1_1,
    matrix_c_1_tile_v_1_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] a_tile_v_26_1 = rf_a_tile_v_1_MPORT_26_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] a_tile_v_26_0 = rf_a_tile_v_0_MPORT_26_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_a_1_T_1 = {a_tile_v_26_1,a_tile_v_26_0,128'h0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 229:35]
  wire [63:0] matrix_b_1_tile_v_2_3 = rf_matrix_b_1_tile_v_3_MPORT_2_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_1_tile_v_2_2 = rf_matrix_b_1_tile_v_2_MPORT_2_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_1_tile_v_2_1 = rf_matrix_b_1_tile_v_1_MPORT_2_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_1_tile_v_2_0 = rf_matrix_b_1_tile_v_0_MPORT_2_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_b_1_T_2 = {matrix_b_1_tile_v_2_3,matrix_b_1_tile_v_2_2,matrix_b_1_tile_v_2_1,
    matrix_b_1_tile_v_2_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] matrix_c_1_tile_v_2_3 = rf_matrix_c_1_tile_v_3_MPORT_2_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_1_tile_v_2_2 = rf_matrix_c_1_tile_v_2_MPORT_2_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_1_tile_v_2_1 = rf_matrix_c_1_tile_v_1_MPORT_2_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_1_tile_v_2_0 = rf_matrix_c_1_tile_v_0_MPORT_2_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_c_1_T_2 = {matrix_c_1_tile_v_2_3,matrix_c_1_tile_v_2_2,matrix_c_1_tile_v_2_1,
    matrix_c_1_tile_v_2_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] a_tile_v_27_3 = rf_a_tile_v_3_MPORT_9_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] a_tile_v_27_2 = rf_a_tile_v_2_MPORT_9_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] a_tile_v_27_1 = rf_a_tile_v_1_MPORT_27_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] a_tile_v_27_0 = rf_a_tile_v_0_MPORT_27_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] a_27 = {a_tile_v_27_3,a_tile_v_27_2,a_tile_v_27_1,a_tile_v_27_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] matrix_b_1_tile_v_3_3 = rf_matrix_b_1_tile_v_3_MPORT_3_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_1_tile_v_3_2 = rf_matrix_b_1_tile_v_2_MPORT_3_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_1_tile_v_3_1 = rf_matrix_b_1_tile_v_1_MPORT_3_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_1_tile_v_3_0 = rf_matrix_b_1_tile_v_0_MPORT_3_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_b_1_T_3 = {matrix_b_1_tile_v_3_3,matrix_b_1_tile_v_3_2,matrix_b_1_tile_v_3_1,
    matrix_b_1_tile_v_3_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] matrix_c_1_tile_v_3_3 = rf_matrix_c_1_tile_v_3_MPORT_3_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_1_tile_v_3_2 = rf_matrix_c_1_tile_v_2_MPORT_3_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_1_tile_v_3_1 = rf_matrix_c_1_tile_v_1_MPORT_3_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_1_tile_v_3_0 = rf_matrix_c_1_tile_v_0_MPORT_3_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_c_1_T_3 = {matrix_c_1_tile_v_3_3,matrix_c_1_tile_v_3_2,matrix_c_1_tile_v_3_1,
    matrix_c_1_tile_v_3_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [255:0] _GEN_1600 = io_mixPc ? _matrix_a_1_T_1 : a_27; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 227:30 229:29 234:29]
  wire [255:0] _GEN_1601 = io_mixPc ? _matrix_b_1_T_2 : _matrix_b_1_T_3; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 227:30 230:29 235:29]
  wire [255:0] _GEN_1606 = io_mixPc ? _matrix_c_1_T_2 : _matrix_c_1_T_3; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 227:30 231:29 236:29]
  wire [63:0] a_tile_v_28_1 = rf_a_tile_v_1_MPORT_28_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] a_tile_v_28_0 = rf_a_tile_v_0_MPORT_28_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_a_1_T_2 = {a_tile_v_28_1,a_tile_v_28_0,128'h0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 241:33]
  wire [63:0] matrix_b_1_tile_v_4_3 = rf_matrix_b_1_tile_v_3_MPORT_4_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_1_tile_v_4_2 = rf_matrix_b_1_tile_v_2_MPORT_4_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_1_tile_v_4_1 = rf_matrix_b_1_tile_v_1_MPORT_4_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_1_tile_v_4_0 = rf_matrix_b_1_tile_v_0_MPORT_4_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_b_1_T_4 = {matrix_b_1_tile_v_4_3,matrix_b_1_tile_v_4_2,matrix_b_1_tile_v_4_1,
    matrix_b_1_tile_v_4_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] matrix_c_1_tile_v_4_3 = rf_matrix_c_1_tile_v_3_MPORT_4_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_1_tile_v_4_2 = rf_matrix_c_1_tile_v_2_MPORT_4_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_1_tile_v_4_1 = rf_matrix_c_1_tile_v_1_MPORT_4_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_1_tile_v_4_0 = rf_matrix_c_1_tile_v_0_MPORT_4_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_c_1_T_4 = {matrix_c_1_tile_v_4_3,matrix_c_1_tile_v_4_2,matrix_c_1_tile_v_4_1,
    matrix_c_1_tile_v_4_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] a_tile_v_29_1 = rf_a_tile_v_1_MPORT_29_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] a_tile_v_29_0 = rf_a_tile_v_0_MPORT_29_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_a_1_T_3 = {a_tile_v_29_1,a_tile_v_29_0,128'h0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 247:33]
  wire [63:0] matrix_b_1_tile_v_5_3 = rf_matrix_b_1_tile_v_3_MPORT_5_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_1_tile_v_5_2 = rf_matrix_b_1_tile_v_2_MPORT_5_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_1_tile_v_5_1 = rf_matrix_b_1_tile_v_1_MPORT_5_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_1_tile_v_5_0 = rf_matrix_b_1_tile_v_0_MPORT_5_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_b_1_T_5 = {matrix_b_1_tile_v_5_3,matrix_b_1_tile_v_5_2,matrix_b_1_tile_v_5_1,
    matrix_b_1_tile_v_5_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] matrix_c_1_tile_v_5_3 = rf_matrix_c_1_tile_v_3_MPORT_5_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_1_tile_v_5_2 = rf_matrix_c_1_tile_v_2_MPORT_5_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_1_tile_v_5_1 = rf_matrix_c_1_tile_v_1_MPORT_5_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_1_tile_v_5_0 = rf_matrix_c_1_tile_v_0_MPORT_5_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_c_1_T_5 = {matrix_c_1_tile_v_5_3,matrix_c_1_tile_v_5_2,matrix_c_1_tile_v_5_1,
    matrix_c_1_tile_v_5_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [255:0] _GEN_1615 = 2'h3 == step ? _matrix_a_1_T_3 : matrix_a_1; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 159:21 212:23 247:27]
  wire [255:0] _GEN_1620 = 2'h3 == step ? _matrix_b_1_T_5 : matrix_b_1; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 160:21 212:23 248:27]
  wire [255:0] _GEN_1625 = 2'h3 == step ? _matrix_c_1_T_5 : matrix_c_1; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 161:21 212:23 249:27]
  wire [255:0] _GEN_1630 = 2'h2 == step ? _matrix_a_1_T_2 : _GEN_1615; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 212:23 241:27]
  wire [255:0] _GEN_1635 = 2'h2 == step ? _matrix_b_1_T_4 : _GEN_1620; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 212:23 242:27]
  wire [255:0] _GEN_1640 = 2'h2 == step ? _matrix_c_1_T_4 : _GEN_1625; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 212:23 243:27]
  wire [63:0] a_tile_v_30_1 = rf_a_tile_v_1_MPORT_30_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] a_tile_v_30_0 = rf_a_tile_v_0_MPORT_30_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_a_1_T_4 = {a_tile_v_30_1,a_tile_v_30_0,128'h0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 258:35]
  wire [63:0] matrix_b_1_tile_v_6_3 = rf_matrix_b_1_tile_v_3_MPORT_6_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_1_tile_v_6_2 = rf_matrix_b_1_tile_v_2_MPORT_6_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_1_tile_v_6_1 = rf_matrix_b_1_tile_v_1_MPORT_6_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_1_tile_v_6_0 = rf_matrix_b_1_tile_v_0_MPORT_6_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_b_1_T_6 = {matrix_b_1_tile_v_6_3,matrix_b_1_tile_v_6_2,matrix_b_1_tile_v_6_1,
    matrix_b_1_tile_v_6_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] matrix_c_1_tile_v_6_3 = rf_matrix_c_1_tile_v_3_MPORT_6_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_1_tile_v_6_2 = rf_matrix_c_1_tile_v_2_MPORT_6_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_1_tile_v_6_1 = rf_matrix_c_1_tile_v_1_MPORT_6_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_1_tile_v_6_0 = rf_matrix_c_1_tile_v_0_MPORT_6_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_c_1_T_6 = {matrix_c_1_tile_v_6_3,matrix_c_1_tile_v_6_2,matrix_c_1_tile_v_6_1,
    matrix_c_1_tile_v_6_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] a_tile_v_31_3 = rf_a_tile_v_3_MPORT_10_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] a_tile_v_31_2 = rf_a_tile_v_2_MPORT_10_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] a_tile_v_31_1 = rf_a_tile_v_1_MPORT_31_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] a_tile_v_31_0 = rf_a_tile_v_0_MPORT_31_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] a_31 = {a_tile_v_31_3,a_tile_v_31_2,a_tile_v_31_1,a_tile_v_31_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] matrix_b_1_tile_v_7_3 = rf_matrix_b_1_tile_v_3_MPORT_7_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_1_tile_v_7_2 = rf_matrix_b_1_tile_v_2_MPORT_7_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_1_tile_v_7_1 = rf_matrix_b_1_tile_v_1_MPORT_7_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_1_tile_v_7_0 = rf_matrix_b_1_tile_v_0_MPORT_7_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_b_1_T_7 = {matrix_b_1_tile_v_7_3,matrix_b_1_tile_v_7_2,matrix_b_1_tile_v_7_1,
    matrix_b_1_tile_v_7_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] matrix_c_1_tile_v_7_3 = rf_matrix_c_1_tile_v_3_MPORT_7_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_1_tile_v_7_2 = rf_matrix_c_1_tile_v_2_MPORT_7_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_1_tile_v_7_1 = rf_matrix_c_1_tile_v_1_MPORT_7_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_1_tile_v_7_0 = rf_matrix_c_1_tile_v_0_MPORT_7_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_c_1_T_7 = {matrix_c_1_tile_v_7_3,matrix_c_1_tile_v_7_2,matrix_c_1_tile_v_7_1,
    matrix_c_1_tile_v_7_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [255:0] _GEN_1787 = io_mixPc ? _matrix_a_1_T_4 : a_31; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 256:30 258:29 263:29]
  wire [255:0] _GEN_1788 = io_mixPc ? _matrix_b_1_T_6 : _matrix_b_1_T_7; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 256:30 259:29 264:29]
  wire [255:0] _GEN_1789 = io_mixPc ? _matrix_c_1_T_6 : _matrix_c_1_T_7; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 256:30 260:29 265:29]
  wire [63:0] a_tile_v_32_1 = rf_a_tile_v_1_MPORT_32_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] a_tile_v_32_0 = rf_a_tile_v_0_MPORT_32_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_a_1_T_5 = {a_tile_v_32_1,a_tile_v_32_0,128'h0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 271:35]
  wire [63:0] matrix_b_1_tile_v_8_3 = rf_matrix_b_1_tile_v_3_MPORT_8_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_1_tile_v_8_2 = rf_matrix_b_1_tile_v_2_MPORT_8_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_1_tile_v_8_1 = rf_matrix_b_1_tile_v_1_MPORT_8_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_1_tile_v_8_0 = rf_matrix_b_1_tile_v_0_MPORT_8_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_b_1_T_8 = {matrix_b_1_tile_v_8_3,matrix_b_1_tile_v_8_2,matrix_b_1_tile_v_8_1,
    matrix_b_1_tile_v_8_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] matrix_c_1_tile_v_8_3 = rf_matrix_c_1_tile_v_3_MPORT_8_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_1_tile_v_8_2 = rf_matrix_c_1_tile_v_2_MPORT_8_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_1_tile_v_8_1 = rf_matrix_c_1_tile_v_1_MPORT_8_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_1_tile_v_8_0 = rf_matrix_c_1_tile_v_0_MPORT_8_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_c_1_T_8 = {matrix_c_1_tile_v_8_3,matrix_c_1_tile_v_8_2,matrix_c_1_tile_v_8_1,
    matrix_c_1_tile_v_8_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] a_tile_v_33_3 = rf_a_tile_v_3_MPORT_11_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] a_tile_v_33_2 = rf_a_tile_v_2_MPORT_11_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] a_tile_v_33_1 = rf_a_tile_v_1_MPORT_33_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] a_tile_v_33_0 = rf_a_tile_v_0_MPORT_33_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] a_33 = {a_tile_v_33_3,a_tile_v_33_2,a_tile_v_33_1,a_tile_v_33_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] matrix_b_1_tile_v_9_3 = rf_matrix_b_1_tile_v_3_MPORT_9_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_1_tile_v_9_2 = rf_matrix_b_1_tile_v_2_MPORT_9_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_1_tile_v_9_1 = rf_matrix_b_1_tile_v_1_MPORT_9_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_1_tile_v_9_0 = rf_matrix_b_1_tile_v_0_MPORT_9_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_b_1_T_9 = {matrix_b_1_tile_v_9_3,matrix_b_1_tile_v_9_2,matrix_b_1_tile_v_9_1,
    matrix_b_1_tile_v_9_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] matrix_c_1_tile_v_9_3 = rf_matrix_c_1_tile_v_3_MPORT_9_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_1_tile_v_9_2 = rf_matrix_c_1_tile_v_2_MPORT_9_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_1_tile_v_9_1 = rf_matrix_c_1_tile_v_1_MPORT_9_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_1_tile_v_9_0 = rf_matrix_c_1_tile_v_0_MPORT_9_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_c_1_T_9 = {matrix_c_1_tile_v_9_3,matrix_c_1_tile_v_9_2,matrix_c_1_tile_v_9_1,
    matrix_c_1_tile_v_9_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [255:0] _GEN_1796 = io_mixPc ? _matrix_a_1_T_5 : a_33; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 269:30 271:29 276:29]
  wire [255:0] _GEN_1797 = io_mixPc ? _matrix_b_1_T_8 : _matrix_b_1_T_9; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 269:30 272:29 277:29]
  wire [255:0] _GEN_1798 = io_mixPc ? _matrix_c_1_T_8 : _matrix_c_1_T_9; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 269:30 273:29 278:29]
  wire [63:0] a_tile_v_34_1 = rf_a_tile_v_1_MPORT_34_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] a_tile_v_34_0 = rf_a_tile_v_0_MPORT_34_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_a_1_T_6 = {a_tile_v_34_1,a_tile_v_34_0,128'h0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 283:33]
  wire [63:0] matrix_b_1_tile_v_10_3 = rf_matrix_b_1_tile_v_3_MPORT_10_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_1_tile_v_10_2 = rf_matrix_b_1_tile_v_2_MPORT_10_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_1_tile_v_10_1 = rf_matrix_b_1_tile_v_1_MPORT_10_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_1_tile_v_10_0 = rf_matrix_b_1_tile_v_0_MPORT_10_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_b_1_T_10 = {matrix_b_1_tile_v_10_3,matrix_b_1_tile_v_10_2,matrix_b_1_tile_v_10_1,
    matrix_b_1_tile_v_10_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] matrix_c_1_tile_v_10_3 = rf_matrix_c_1_tile_v_3_MPORT_10_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_1_tile_v_10_2 = rf_matrix_c_1_tile_v_2_MPORT_10_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_1_tile_v_10_1 = rf_matrix_c_1_tile_v_1_MPORT_10_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_1_tile_v_10_0 = rf_matrix_c_1_tile_v_0_MPORT_10_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_c_1_T_10 = {matrix_c_1_tile_v_10_3,matrix_c_1_tile_v_10_2,matrix_c_1_tile_v_10_1,
    matrix_c_1_tile_v_10_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] a_tile_v_35_1 = rf_a_tile_v_1_MPORT_35_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] a_tile_v_35_0 = rf_a_tile_v_0_MPORT_35_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_a_1_T_7 = {a_tile_v_35_1,a_tile_v_35_0,128'h0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 289:33]
  wire [63:0] matrix_b_1_tile_v_11_3 = rf_matrix_b_1_tile_v_3_MPORT_11_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_1_tile_v_11_2 = rf_matrix_b_1_tile_v_2_MPORT_11_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_1_tile_v_11_1 = rf_matrix_b_1_tile_v_1_MPORT_11_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_1_tile_v_11_0 = rf_matrix_b_1_tile_v_0_MPORT_11_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_b_1_T_11 = {matrix_b_1_tile_v_11_3,matrix_b_1_tile_v_11_2,matrix_b_1_tile_v_11_1,
    matrix_b_1_tile_v_11_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] matrix_c_1_tile_v_11_3 = rf_matrix_c_1_tile_v_3_MPORT_11_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_1_tile_v_11_2 = rf_matrix_c_1_tile_v_2_MPORT_11_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_1_tile_v_11_1 = rf_matrix_c_1_tile_v_1_MPORT_11_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_1_tile_v_11_0 = rf_matrix_c_1_tile_v_0_MPORT_11_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_c_1_T_11 = {matrix_c_1_tile_v_11_3,matrix_c_1_tile_v_11_2,matrix_c_1_tile_v_11_1,
    matrix_c_1_tile_v_11_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [255:0] _GEN_1803 = _T_4 ? _matrix_a_1_T_7 : matrix_a_1; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 159:21 254:24 289:27]
  wire [255:0] _GEN_1808 = _T_4 ? _matrix_b_1_T_11 : matrix_b_1; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 160:21 254:24 290:27]
  wire [255:0] _GEN_1813 = _T_4 ? _matrix_c_1_T_11 : matrix_c_1; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 161:21 254:24 291:27]
  wire [255:0] _GEN_1818 = _T_3 ? _matrix_a_1_T_6 : _GEN_1803; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 254:24 283:27]
  wire [255:0] _GEN_1823 = _T_3 ? _matrix_b_1_T_10 : _GEN_1808; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 254:24 284:27]
  wire [255:0] _GEN_1828 = _T_3 ? _matrix_c_1_T_10 : _GEN_1813; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 254:24 285:27]
  wire [255:0] _GEN_1845 = _T_2 ? _GEN_1796 : _GEN_1818; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 254:24]
  wire [255:0] _GEN_1850 = _T_2 ? _GEN_1797 : _GEN_1823; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 254:24]
  wire [255:0] _GEN_1855 = _T_2 ? _GEN_1798 : _GEN_1828; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 254:24]
  wire [63:0] a_tile_v_36_1 = rf_a_tile_v_1_MPORT_36_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] a_tile_v_36_0 = rf_a_tile_v_0_MPORT_36_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_a_1_T_8 = {a_tile_v_36_1,a_tile_v_36_0,128'h0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 300:35]
  wire [63:0] matrix_b_1_tile_v_12_3 = rf_matrix_b_1_tile_v_3_MPORT_12_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_1_tile_v_12_2 = rf_matrix_b_1_tile_v_2_MPORT_12_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_1_tile_v_12_1 = rf_matrix_b_1_tile_v_1_MPORT_12_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_1_tile_v_12_0 = rf_matrix_b_1_tile_v_0_MPORT_12_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_b_1_T_12 = {matrix_b_1_tile_v_12_3,matrix_b_1_tile_v_12_2,matrix_b_1_tile_v_12_1,
    matrix_b_1_tile_v_12_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] matrix_c_1_tile_v_12_3 = rf_matrix_c_1_tile_v_3_MPORT_12_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_1_tile_v_12_2 = rf_matrix_c_1_tile_v_2_MPORT_12_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_1_tile_v_12_1 = rf_matrix_c_1_tile_v_1_MPORT_12_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_1_tile_v_12_0 = rf_matrix_c_1_tile_v_0_MPORT_12_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_c_1_T_12 = {matrix_c_1_tile_v_12_3,matrix_c_1_tile_v_12_2,matrix_c_1_tile_v_12_1,
    matrix_c_1_tile_v_12_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] a_tile_v_37_3 = rf_a_tile_v_3_MPORT_12_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] a_tile_v_37_2 = rf_a_tile_v_2_MPORT_12_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] a_tile_v_37_1 = rf_a_tile_v_1_MPORT_37_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] a_tile_v_37_0 = rf_a_tile_v_0_MPORT_37_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] a_37 = {a_tile_v_37_3,a_tile_v_37_2,a_tile_v_37_1,a_tile_v_37_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] matrix_b_1_tile_v_13_3 = rf_matrix_b_1_tile_v_3_MPORT_13_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_1_tile_v_13_2 = rf_matrix_b_1_tile_v_2_MPORT_13_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_1_tile_v_13_1 = rf_matrix_b_1_tile_v_1_MPORT_13_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_1_tile_v_13_0 = rf_matrix_b_1_tile_v_0_MPORT_13_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_b_1_T_13 = {matrix_b_1_tile_v_13_3,matrix_b_1_tile_v_13_2,matrix_b_1_tile_v_13_1,
    matrix_b_1_tile_v_13_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] matrix_c_1_tile_v_13_3 = rf_matrix_c_1_tile_v_3_MPORT_13_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_1_tile_v_13_2 = rf_matrix_c_1_tile_v_2_MPORT_13_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_1_tile_v_13_1 = rf_matrix_c_1_tile_v_1_MPORT_13_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_1_tile_v_13_0 = rf_matrix_c_1_tile_v_0_MPORT_13_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_c_1_T_13 = {matrix_c_1_tile_v_13_3,matrix_c_1_tile_v_13_2,matrix_c_1_tile_v_13_1,
    matrix_c_1_tile_v_13_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [255:0] _GEN_1975 = io_mixPc ? _matrix_a_1_T_8 : a_37; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 298:30 300:29 305:29]
  wire [255:0] _GEN_1976 = io_mixPc ? _matrix_b_1_T_12 : _matrix_b_1_T_13; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 298:30 301:29 306:29]
  wire [255:0] _GEN_1977 = io_mixPc ? _matrix_c_1_T_12 : _matrix_c_1_T_13; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 298:30 302:29 307:29]
  wire [63:0] a_tile_v_38_1 = rf_a_tile_v_1_MPORT_38_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] a_tile_v_38_0 = rf_a_tile_v_0_MPORT_38_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_a_1_T_9 = {a_tile_v_38_1,a_tile_v_38_0,128'h0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 313:35]
  wire [63:0] matrix_b_1_tile_v_14_3 = rf_matrix_b_1_tile_v_3_MPORT_14_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_1_tile_v_14_2 = rf_matrix_b_1_tile_v_2_MPORT_14_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_1_tile_v_14_1 = rf_matrix_b_1_tile_v_1_MPORT_14_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_1_tile_v_14_0 = rf_matrix_b_1_tile_v_0_MPORT_14_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_b_1_T_14 = {matrix_b_1_tile_v_14_3,matrix_b_1_tile_v_14_2,matrix_b_1_tile_v_14_1,
    matrix_b_1_tile_v_14_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] matrix_c_1_tile_v_14_3 = rf_matrix_c_1_tile_v_3_MPORT_14_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_1_tile_v_14_2 = rf_matrix_c_1_tile_v_2_MPORT_14_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_1_tile_v_14_1 = rf_matrix_c_1_tile_v_1_MPORT_14_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_1_tile_v_14_0 = rf_matrix_c_1_tile_v_0_MPORT_14_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_c_1_T_14 = {matrix_c_1_tile_v_14_3,matrix_c_1_tile_v_14_2,matrix_c_1_tile_v_14_1,
    matrix_c_1_tile_v_14_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] a_tile_v_39_3 = rf_a_tile_v_3_MPORT_13_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] a_tile_v_39_2 = rf_a_tile_v_2_MPORT_13_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] a_tile_v_39_1 = rf_a_tile_v_1_MPORT_39_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] a_tile_v_39_0 = rf_a_tile_v_0_MPORT_39_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] a_39 = {a_tile_v_39_3,a_tile_v_39_2,a_tile_v_39_1,a_tile_v_39_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] matrix_b_1_tile_v_15_3 = rf_matrix_b_1_tile_v_3_MPORT_15_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_1_tile_v_15_2 = rf_matrix_b_1_tile_v_2_MPORT_15_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_1_tile_v_15_1 = rf_matrix_b_1_tile_v_1_MPORT_15_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_1_tile_v_15_0 = rf_matrix_b_1_tile_v_0_MPORT_15_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_b_1_T_15 = {matrix_b_1_tile_v_15_3,matrix_b_1_tile_v_15_2,matrix_b_1_tile_v_15_1,
    matrix_b_1_tile_v_15_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] matrix_c_1_tile_v_15_3 = rf_matrix_c_1_tile_v_3_MPORT_15_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_1_tile_v_15_2 = rf_matrix_c_1_tile_v_2_MPORT_15_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_1_tile_v_15_1 = rf_matrix_c_1_tile_v_1_MPORT_15_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_1_tile_v_15_0 = rf_matrix_c_1_tile_v_0_MPORT_15_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_c_1_T_15 = {matrix_c_1_tile_v_15_3,matrix_c_1_tile_v_15_2,matrix_c_1_tile_v_15_1,
    matrix_c_1_tile_v_15_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [255:0] _GEN_1984 = io_mixPc ? _matrix_a_1_T_9 : a_39; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 311:30 313:29 318:29]
  wire [255:0] _GEN_1985 = io_mixPc ? _matrix_b_1_T_14 : _matrix_b_1_T_15; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 311:30 314:29 319:29]
  wire [255:0] _GEN_1986 = io_mixPc ? _matrix_c_1_T_14 : _matrix_c_1_T_15; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 311:30 315:29 320:29]
  wire [63:0] a_tile_v_40_1 = rf_a_tile_v_1_MPORT_40_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] a_tile_v_40_0 = rf_a_tile_v_0_MPORT_40_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_a_1_T_10 = {a_tile_v_40_1,a_tile_v_40_0,128'h0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 325:33]
  wire [63:0] matrix_b_1_tile_v_16_3 = rf_matrix_b_1_tile_v_3_MPORT_16_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_1_tile_v_16_2 = rf_matrix_b_1_tile_v_2_MPORT_16_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_1_tile_v_16_1 = rf_matrix_b_1_tile_v_1_MPORT_16_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_1_tile_v_16_0 = rf_matrix_b_1_tile_v_0_MPORT_16_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_b_1_T_16 = {matrix_b_1_tile_v_16_3,matrix_b_1_tile_v_16_2,matrix_b_1_tile_v_16_1,
    matrix_b_1_tile_v_16_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] matrix_c_1_tile_v_16_3 = rf_matrix_c_1_tile_v_3_MPORT_16_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_1_tile_v_16_2 = rf_matrix_c_1_tile_v_2_MPORT_16_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_1_tile_v_16_1 = rf_matrix_c_1_tile_v_1_MPORT_16_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_1_tile_v_16_0 = rf_matrix_c_1_tile_v_0_MPORT_16_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_c_1_T_16 = {matrix_c_1_tile_v_16_3,matrix_c_1_tile_v_16_2,matrix_c_1_tile_v_16_1,
    matrix_c_1_tile_v_16_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] a_tile_v_41_1 = rf_a_tile_v_1_MPORT_41_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] a_tile_v_41_0 = rf_a_tile_v_0_MPORT_41_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_a_1_T_11 = {a_tile_v_41_1,a_tile_v_41_0,128'h0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 331:33]
  wire [63:0] matrix_b_1_tile_v_17_3 = rf_matrix_b_1_tile_v_3_MPORT_17_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_1_tile_v_17_2 = rf_matrix_b_1_tile_v_2_MPORT_17_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_1_tile_v_17_1 = rf_matrix_b_1_tile_v_1_MPORT_17_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_1_tile_v_17_0 = rf_matrix_b_1_tile_v_0_MPORT_17_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_b_1_T_17 = {matrix_b_1_tile_v_17_3,matrix_b_1_tile_v_17_2,matrix_b_1_tile_v_17_1,
    matrix_b_1_tile_v_17_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] matrix_c_1_tile_v_17_3 = rf_matrix_c_1_tile_v_3_MPORT_17_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_1_tile_v_17_2 = rf_matrix_c_1_tile_v_2_MPORT_17_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_1_tile_v_17_1 = rf_matrix_c_1_tile_v_1_MPORT_17_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_1_tile_v_17_0 = rf_matrix_c_1_tile_v_0_MPORT_17_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_c_1_T_17 = {matrix_c_1_tile_v_17_3,matrix_c_1_tile_v_17_2,matrix_c_1_tile_v_17_1,
    matrix_c_1_tile_v_17_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [255:0] _GEN_1991 = _T_4 ? _matrix_a_1_T_11 : matrix_a_1; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 159:21 296:24 331:27]
  wire [255:0] _GEN_1996 = _T_4 ? _matrix_b_1_T_17 : matrix_b_1; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 160:21 296:24 332:27]
  wire [255:0] _GEN_2001 = _T_4 ? _matrix_c_1_T_17 : matrix_c_1; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 161:21 296:24 333:27]
  wire [255:0] _GEN_2006 = _T_3 ? _matrix_a_1_T_10 : _GEN_1991; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 296:24 325:27]
  wire [255:0] _GEN_2011 = _T_3 ? _matrix_b_1_T_16 : _GEN_1996; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 296:24 326:27]
  wire [255:0] _GEN_2016 = _T_3 ? _matrix_c_1_T_16 : _GEN_2001; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 296:24 327:27]
  wire [255:0] _GEN_2033 = _T_2 ? _GEN_1984 : _GEN_2006; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 296:24]
  wire [255:0] _GEN_2038 = _T_2 ? _GEN_1985 : _GEN_2011; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 296:24]
  wire [255:0] _GEN_2043 = _T_2 ? _GEN_1986 : _GEN_2016; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 296:24]
  wire [255:0] _GEN_2086 = _T_1 ? _GEN_1975 : _GEN_2033; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 296:24]
  wire [255:0] _GEN_2091 = _T_1 ? _GEN_1976 : _GEN_2038; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 296:24]
  wire [255:0] _GEN_2096 = _T_1 ? _GEN_1977 : _GEN_2043; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 296:24]
  wire [63:0] a_tile_v_42_1 = rf_a_tile_v_1_MPORT_42_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] a_tile_v_42_0 = rf_a_tile_v_0_MPORT_42_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_a_1_T_12 = {a_tile_v_42_1,a_tile_v_42_0,128'h0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 342:35]
  wire [63:0] matrix_b_1_tile_v_18_3 = rf_matrix_b_1_tile_v_3_MPORT_18_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_1_tile_v_18_2 = rf_matrix_b_1_tile_v_2_MPORT_18_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_1_tile_v_18_1 = rf_matrix_b_1_tile_v_1_MPORT_18_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_1_tile_v_18_0 = rf_matrix_b_1_tile_v_0_MPORT_18_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_b_1_T_18 = {matrix_b_1_tile_v_18_3,matrix_b_1_tile_v_18_2,matrix_b_1_tile_v_18_1,
    matrix_b_1_tile_v_18_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] matrix_c_1_tile_v_18_3 = rf_matrix_c_1_tile_v_3_MPORT_18_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_1_tile_v_18_2 = rf_matrix_c_1_tile_v_2_MPORT_18_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_1_tile_v_18_1 = rf_matrix_c_1_tile_v_1_MPORT_18_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_1_tile_v_18_0 = rf_matrix_c_1_tile_v_0_MPORT_18_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_c_1_T_18 = {matrix_c_1_tile_v_18_3,matrix_c_1_tile_v_18_2,matrix_c_1_tile_v_18_1,
    matrix_c_1_tile_v_18_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] a_tile_v_43_3 = rf_a_tile_v_3_MPORT_14_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] a_tile_v_43_2 = rf_a_tile_v_2_MPORT_14_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] a_tile_v_43_1 = rf_a_tile_v_1_MPORT_43_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] a_tile_v_43_0 = rf_a_tile_v_0_MPORT_43_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] a_43 = {a_tile_v_43_3,a_tile_v_43_2,a_tile_v_43_1,a_tile_v_43_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] matrix_b_1_tile_v_19_3 = rf_matrix_b_1_tile_v_3_MPORT_19_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_1_tile_v_19_2 = rf_matrix_b_1_tile_v_2_MPORT_19_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_1_tile_v_19_1 = rf_matrix_b_1_tile_v_1_MPORT_19_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_1_tile_v_19_0 = rf_matrix_b_1_tile_v_0_MPORT_19_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_b_1_T_19 = {matrix_b_1_tile_v_19_3,matrix_b_1_tile_v_19_2,matrix_b_1_tile_v_19_1,
    matrix_b_1_tile_v_19_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] matrix_c_1_tile_v_19_3 = rf_matrix_c_1_tile_v_3_MPORT_19_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_1_tile_v_19_2 = rf_matrix_c_1_tile_v_2_MPORT_19_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_1_tile_v_19_1 = rf_matrix_c_1_tile_v_1_MPORT_19_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_1_tile_v_19_0 = rf_matrix_c_1_tile_v_0_MPORT_19_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_c_1_T_19 = {matrix_c_1_tile_v_19_3,matrix_c_1_tile_v_19_2,matrix_c_1_tile_v_19_1,
    matrix_c_1_tile_v_19_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [255:0] _GEN_2163 = io_mixPc ? _matrix_a_1_T_12 : a_43; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 340:30 342:29 347:29]
  wire [255:0] _GEN_2164 = io_mixPc ? _matrix_b_1_T_18 : _matrix_b_1_T_19; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 340:30 343:29 348:29]
  wire [255:0] _GEN_2165 = io_mixPc ? _matrix_c_1_T_18 : _matrix_c_1_T_19; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 340:30 344:29 349:29]
  wire [63:0] a_tile_v_44_1 = rf_a_tile_v_1_MPORT_44_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] a_tile_v_44_0 = rf_a_tile_v_0_MPORT_44_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_a_1_T_13 = {a_tile_v_44_1,a_tile_v_44_0,128'h0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 355:35]
  wire [63:0] matrix_b_1_tile_v_20_3 = rf_matrix_b_1_tile_v_3_MPORT_20_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_1_tile_v_20_2 = rf_matrix_b_1_tile_v_2_MPORT_20_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_1_tile_v_20_1 = rf_matrix_b_1_tile_v_1_MPORT_20_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_1_tile_v_20_0 = rf_matrix_b_1_tile_v_0_MPORT_20_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_b_1_T_20 = {matrix_b_1_tile_v_20_3,matrix_b_1_tile_v_20_2,matrix_b_1_tile_v_20_1,
    matrix_b_1_tile_v_20_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] matrix_c_1_tile_v_20_3 = rf_matrix_c_1_tile_v_3_MPORT_20_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_1_tile_v_20_2 = rf_matrix_c_1_tile_v_2_MPORT_20_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_1_tile_v_20_1 = rf_matrix_c_1_tile_v_1_MPORT_20_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_1_tile_v_20_0 = rf_matrix_c_1_tile_v_0_MPORT_20_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_c_1_T_20 = {matrix_c_1_tile_v_20_3,matrix_c_1_tile_v_20_2,matrix_c_1_tile_v_20_1,
    matrix_c_1_tile_v_20_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] a_tile_v_45_3 = rf_a_tile_v_3_MPORT_15_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] a_tile_v_45_2 = rf_a_tile_v_2_MPORT_15_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] a_tile_v_45_1 = rf_a_tile_v_1_MPORT_45_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] a_tile_v_45_0 = rf_a_tile_v_0_MPORT_45_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] a_45 = {a_tile_v_45_3,a_tile_v_45_2,a_tile_v_45_1,a_tile_v_45_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] matrix_b_1_tile_v_21_3 = rf_matrix_b_1_tile_v_3_MPORT_21_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_1_tile_v_21_2 = rf_matrix_b_1_tile_v_2_MPORT_21_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_1_tile_v_21_1 = rf_matrix_b_1_tile_v_1_MPORT_21_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_1_tile_v_21_0 = rf_matrix_b_1_tile_v_0_MPORT_21_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_b_1_T_21 = {matrix_b_1_tile_v_21_3,matrix_b_1_tile_v_21_2,matrix_b_1_tile_v_21_1,
    matrix_b_1_tile_v_21_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] matrix_c_1_tile_v_21_3 = rf_matrix_c_1_tile_v_3_MPORT_21_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_1_tile_v_21_2 = rf_matrix_c_1_tile_v_2_MPORT_21_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_1_tile_v_21_1 = rf_matrix_c_1_tile_v_1_MPORT_21_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_1_tile_v_21_0 = rf_matrix_c_1_tile_v_0_MPORT_21_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_c_1_T_21 = {matrix_c_1_tile_v_21_3,matrix_c_1_tile_v_21_2,matrix_c_1_tile_v_21_1,
    matrix_c_1_tile_v_21_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [255:0] _GEN_2172 = io_mixPc ? _matrix_a_1_T_13 : a_45; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 353:30 355:29 360:29]
  wire [255:0] _GEN_2173 = io_mixPc ? _matrix_b_1_T_20 : _matrix_b_1_T_21; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 353:30 356:29 361:29]
  wire [255:0] _GEN_2174 = io_mixPc ? _matrix_c_1_T_20 : _matrix_c_1_T_21; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 353:30 357:29 362:29]
  wire [63:0] a_tile_v_46_1 = rf_a_tile_v_1_MPORT_46_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] a_tile_v_46_0 = rf_a_tile_v_0_MPORT_46_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_a_1_T_14 = {a_tile_v_46_1,a_tile_v_46_0,128'h0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 367:33]
  wire [63:0] matrix_b_1_tile_v_22_3 = rf_matrix_b_1_tile_v_3_MPORT_22_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_1_tile_v_22_2 = rf_matrix_b_1_tile_v_2_MPORT_22_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_1_tile_v_22_1 = rf_matrix_b_1_tile_v_1_MPORT_22_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_1_tile_v_22_0 = rf_matrix_b_1_tile_v_0_MPORT_22_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_b_1_T_22 = {matrix_b_1_tile_v_22_3,matrix_b_1_tile_v_22_2,matrix_b_1_tile_v_22_1,
    matrix_b_1_tile_v_22_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] matrix_c_1_tile_v_22_3 = rf_matrix_c_1_tile_v_3_MPORT_22_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_1_tile_v_22_2 = rf_matrix_c_1_tile_v_2_MPORT_22_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_1_tile_v_22_1 = rf_matrix_c_1_tile_v_1_MPORT_22_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_1_tile_v_22_0 = rf_matrix_c_1_tile_v_0_MPORT_22_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_c_1_T_22 = {matrix_c_1_tile_v_22_3,matrix_c_1_tile_v_22_2,matrix_c_1_tile_v_22_1,
    matrix_c_1_tile_v_22_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] a_tile_v_47_1 = rf_a_tile_v_1_MPORT_47_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] a_tile_v_47_0 = rf_a_tile_v_0_MPORT_47_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_a_1_T_15 = {a_tile_v_47_1,a_tile_v_47_0,128'h0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 373:33]
  wire [63:0] matrix_b_1_tile_v_23_3 = rf_matrix_b_1_tile_v_3_MPORT_23_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_1_tile_v_23_2 = rf_matrix_b_1_tile_v_2_MPORT_23_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_1_tile_v_23_1 = rf_matrix_b_1_tile_v_1_MPORT_23_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_1_tile_v_23_0 = rf_matrix_b_1_tile_v_0_MPORT_23_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_b_1_T_23 = {matrix_b_1_tile_v_23_3,matrix_b_1_tile_v_23_2,matrix_b_1_tile_v_23_1,
    matrix_b_1_tile_v_23_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] matrix_c_1_tile_v_23_3 = rf_matrix_c_1_tile_v_3_MPORT_23_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_1_tile_v_23_2 = rf_matrix_c_1_tile_v_2_MPORT_23_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_1_tile_v_23_1 = rf_matrix_c_1_tile_v_1_MPORT_23_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_1_tile_v_23_0 = rf_matrix_c_1_tile_v_0_MPORT_23_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_c_1_T_23 = {matrix_c_1_tile_v_23_3,matrix_c_1_tile_v_23_2,matrix_c_1_tile_v_23_1,
    matrix_c_1_tile_v_23_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [255:0] _GEN_2179 = _T_4 ? _matrix_a_1_T_15 : matrix_a_1; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 159:21 338:24 373:27]
  wire [255:0] _GEN_2184 = _T_4 ? _matrix_b_1_T_23 : matrix_b_1; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 160:21 338:24 374:27]
  wire [255:0] _GEN_2189 = _T_4 ? _matrix_c_1_T_23 : matrix_c_1; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 161:21 338:24 375:27]
  wire [255:0] _GEN_2194 = _T_3 ? _matrix_a_1_T_14 : _GEN_2179; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 338:24 367:27]
  wire [255:0] _GEN_2199 = _T_3 ? _matrix_b_1_T_22 : _GEN_2184; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 338:24 368:27]
  wire [255:0] _GEN_2204 = _T_3 ? _matrix_c_1_T_22 : _GEN_2189; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 338:24 369:27]
  wire [255:0] _GEN_2221 = _T_2 ? _GEN_2172 : _GEN_2194; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 338:24]
  wire [255:0] _GEN_2226 = _T_2 ? _GEN_2173 : _GEN_2199; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 338:24]
  wire [255:0] _GEN_2231 = _T_2 ? _GEN_2174 : _GEN_2204; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 338:24]
  wire [255:0] _GEN_2274 = _T_1 ? _GEN_2163 : _GEN_2221; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 338:24]
  wire [255:0] _GEN_2279 = _T_1 ? _GEN_2164 : _GEN_2226; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 338:24]
  wire [255:0] _GEN_2284 = _T_1 ? _GEN_2165 : _GEN_2231; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 338:24]
  wire [255:0] _GEN_2353 = 2'h3 == set ? _GEN_2274 : matrix_a_1; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 210:18 159:21]
  wire [255:0] _GEN_2358 = 2'h3 == set ? _GEN_2279 : matrix_b_1; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 210:18 160:21]
  wire [255:0] _GEN_2363 = 2'h3 == set ? _GEN_2284 : matrix_c_1; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 210:18 161:21]
  wire [63:0] a_tile_v_48_0 = rf_a_tile_v_0_MPORT_48_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_a_2_T = {64'h0,a_tile_v_48_0,128'h0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 216:35]
  wire [63:0] matrix_b_2_tile_v__3 = rf_matrix_b_2_tile_v_3_MPORT_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_2_tile_v__2 = rf_matrix_b_2_tile_v_2_MPORT_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_2_tile_v__1 = rf_matrix_b_2_tile_v_1_MPORT_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_2_tile_v__0 = rf_matrix_b_2_tile_v_0_MPORT_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_b_2_T = {matrix_b_2_tile_v__3,matrix_b_2_tile_v__2,matrix_b_2_tile_v__1,matrix_b_2_tile_v__0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] matrix_c_2_tile_v__3 = rf_matrix_c_2_tile_v_3_MPORT_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_2_tile_v__2 = rf_matrix_c_2_tile_v_2_MPORT_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_2_tile_v__1 = rf_matrix_c_2_tile_v_1_MPORT_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_2_tile_v__0 = rf_matrix_c_2_tile_v_0_MPORT_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_c_2_T = {matrix_c_2_tile_v__3,matrix_c_2_tile_v__2,matrix_c_2_tile_v__1,matrix_c_2_tile_v__0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] a_tile_v_49_2 = rf_a_tile_v_2_MPORT_16_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] a_tile_v_49_1 = rf_a_tile_v_1_MPORT_49_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] a_tile_v_49_0 = rf_a_tile_v_0_MPORT_49_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] a_49 = {64'h0,a_tile_v_49_2,a_tile_v_49_1,a_tile_v_49_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] matrix_b_2_tile_v_1_3 = rf_matrix_b_2_tile_v_3_MPORT_1_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_2_tile_v_1_2 = rf_matrix_b_2_tile_v_2_MPORT_1_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_2_tile_v_1_1 = rf_matrix_b_2_tile_v_1_MPORT_1_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_2_tile_v_1_0 = rf_matrix_b_2_tile_v_0_MPORT_1_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_b_2_T_1 = {matrix_b_2_tile_v_1_3,matrix_b_2_tile_v_1_2,matrix_b_2_tile_v_1_1,
    matrix_b_2_tile_v_1_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] matrix_c_2_tile_v_1_3 = rf_matrix_c_2_tile_v_3_MPORT_1_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_2_tile_v_1_2 = rf_matrix_c_2_tile_v_2_MPORT_1_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_2_tile_v_1_1 = rf_matrix_c_2_tile_v_1_MPORT_1_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_2_tile_v_1_0 = rf_matrix_c_2_tile_v_0_MPORT_1_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_c_2_T_1 = {matrix_c_2_tile_v_1_3,matrix_c_2_tile_v_1_2,matrix_c_2_tile_v_1_1,
    matrix_c_2_tile_v_1_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] a_tile_v_50_1 = rf_a_tile_v_1_MPORT_50_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] a_tile_v_50_0 = rf_a_tile_v_0_MPORT_50_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_a_2_T_1 = {a_tile_v_50_1,a_tile_v_50_0,128'h0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 229:35]
  wire [63:0] matrix_b_2_tile_v_2_3 = rf_matrix_b_2_tile_v_3_MPORT_2_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_2_tile_v_2_2 = rf_matrix_b_2_tile_v_2_MPORT_2_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_2_tile_v_2_1 = rf_matrix_b_2_tile_v_1_MPORT_2_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_2_tile_v_2_0 = rf_matrix_b_2_tile_v_0_MPORT_2_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_b_2_T_2 = {matrix_b_2_tile_v_2_3,matrix_b_2_tile_v_2_2,matrix_b_2_tile_v_2_1,
    matrix_b_2_tile_v_2_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] matrix_c_2_tile_v_2_3 = rf_matrix_c_2_tile_v_3_MPORT_2_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_2_tile_v_2_2 = rf_matrix_c_2_tile_v_2_MPORT_2_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_2_tile_v_2_1 = rf_matrix_c_2_tile_v_1_MPORT_2_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_2_tile_v_2_0 = rf_matrix_c_2_tile_v_0_MPORT_2_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_c_2_T_2 = {matrix_c_2_tile_v_2_3,matrix_c_2_tile_v_2_2,matrix_c_2_tile_v_2_1,
    matrix_c_2_tile_v_2_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] a_tile_v_51_2 = rf_a_tile_v_2_MPORT_17_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] a_tile_v_51_1 = rf_a_tile_v_1_MPORT_51_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] a_tile_v_51_0 = rf_a_tile_v_0_MPORT_51_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] a_51 = {64'h0,a_tile_v_51_2,a_tile_v_51_1,a_tile_v_51_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] matrix_b_2_tile_v_3_3 = rf_matrix_b_2_tile_v_3_MPORT_3_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_2_tile_v_3_2 = rf_matrix_b_2_tile_v_2_MPORT_3_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_2_tile_v_3_1 = rf_matrix_b_2_tile_v_1_MPORT_3_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_2_tile_v_3_0 = rf_matrix_b_2_tile_v_0_MPORT_3_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_b_2_T_3 = {matrix_b_2_tile_v_3_3,matrix_b_2_tile_v_3_2,matrix_b_2_tile_v_3_1,
    matrix_b_2_tile_v_3_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] matrix_c_2_tile_v_3_3 = rf_matrix_c_2_tile_v_3_MPORT_3_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_2_tile_v_3_2 = rf_matrix_c_2_tile_v_2_MPORT_3_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_2_tile_v_3_1 = rf_matrix_c_2_tile_v_1_MPORT_3_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_2_tile_v_3_0 = rf_matrix_c_2_tile_v_0_MPORT_3_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_c_2_T_3 = {matrix_c_2_tile_v_3_3,matrix_c_2_tile_v_3_2,matrix_c_2_tile_v_3_1,
    matrix_c_2_tile_v_3_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [255:0] _GEN_3140 = io_mixPc ? _matrix_a_2_T_1 : a_51; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 227:30 229:29 234:29]
  wire [255:0] _GEN_3141 = io_mixPc ? _matrix_b_2_T_2 : _matrix_b_2_T_3; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 227:30 230:29 235:29]
  wire [255:0] _GEN_3146 = io_mixPc ? _matrix_c_2_T_2 : _matrix_c_2_T_3; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 227:30 231:29 236:29]
  wire [63:0] a_tile_v_52_0 = rf_a_tile_v_0_MPORT_52_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_a_2_T_2 = {64'h0,a_tile_v_52_0,128'h0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 241:33]
  wire [63:0] matrix_b_2_tile_v_4_3 = rf_matrix_b_2_tile_v_3_MPORT_4_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_2_tile_v_4_2 = rf_matrix_b_2_tile_v_2_MPORT_4_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_2_tile_v_4_1 = rf_matrix_b_2_tile_v_1_MPORT_4_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_2_tile_v_4_0 = rf_matrix_b_2_tile_v_0_MPORT_4_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_b_2_T_4 = {matrix_b_2_tile_v_4_3,matrix_b_2_tile_v_4_2,matrix_b_2_tile_v_4_1,
    matrix_b_2_tile_v_4_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] matrix_c_2_tile_v_4_3 = rf_matrix_c_2_tile_v_3_MPORT_4_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_2_tile_v_4_2 = rf_matrix_c_2_tile_v_2_MPORT_4_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_2_tile_v_4_1 = rf_matrix_c_2_tile_v_1_MPORT_4_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_2_tile_v_4_0 = rf_matrix_c_2_tile_v_0_MPORT_4_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_c_2_T_4 = {matrix_c_2_tile_v_4_3,matrix_c_2_tile_v_4_2,matrix_c_2_tile_v_4_1,
    matrix_c_2_tile_v_4_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] a_tile_v_53_1 = rf_a_tile_v_1_MPORT_53_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] a_tile_v_53_0 = rf_a_tile_v_0_MPORT_53_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_a_2_T_3 = {a_tile_v_53_1,a_tile_v_53_0,128'h0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 247:33]
  wire [63:0] matrix_b_2_tile_v_5_3 = rf_matrix_b_2_tile_v_3_MPORT_5_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_2_tile_v_5_2 = rf_matrix_b_2_tile_v_2_MPORT_5_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_2_tile_v_5_1 = rf_matrix_b_2_tile_v_1_MPORT_5_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_2_tile_v_5_0 = rf_matrix_b_2_tile_v_0_MPORT_5_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_b_2_T_5 = {matrix_b_2_tile_v_5_3,matrix_b_2_tile_v_5_2,matrix_b_2_tile_v_5_1,
    matrix_b_2_tile_v_5_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] matrix_c_2_tile_v_5_3 = rf_matrix_c_2_tile_v_3_MPORT_5_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_2_tile_v_5_2 = rf_matrix_c_2_tile_v_2_MPORT_5_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_2_tile_v_5_1 = rf_matrix_c_2_tile_v_1_MPORT_5_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_2_tile_v_5_0 = rf_matrix_c_2_tile_v_0_MPORT_5_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_c_2_T_5 = {matrix_c_2_tile_v_5_3,matrix_c_2_tile_v_5_2,matrix_c_2_tile_v_5_1,
    matrix_c_2_tile_v_5_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [255:0] _GEN_3155 = 2'h3 == step ? _matrix_a_2_T_3 : matrix_a_2; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 159:21 212:23 247:27]
  wire [255:0] _GEN_3160 = 2'h3 == step ? _matrix_b_2_T_5 : matrix_b_2; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 160:21 212:23 248:27]
  wire [255:0] _GEN_3165 = 2'h3 == step ? _matrix_c_2_T_5 : matrix_c_2; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 161:21 212:23 249:27]
  wire [255:0] _GEN_3170 = 2'h2 == step ? _matrix_a_2_T_2 : _GEN_3155; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 212:23 241:27]
  wire [255:0] _GEN_3175 = 2'h2 == step ? _matrix_b_2_T_4 : _GEN_3160; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 212:23 242:27]
  wire [255:0] _GEN_3180 = 2'h2 == step ? _matrix_c_2_T_4 : _GEN_3165; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 212:23 243:27]
  wire [63:0] a_tile_v_54_1 = rf_a_tile_v_1_MPORT_54_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] a_tile_v_54_0 = rf_a_tile_v_0_MPORT_54_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_a_2_T_4 = {a_tile_v_54_1,a_tile_v_54_0,128'h0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 258:35]
  wire [63:0] matrix_b_2_tile_v_6_3 = rf_matrix_b_2_tile_v_3_MPORT_6_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_2_tile_v_6_2 = rf_matrix_b_2_tile_v_2_MPORT_6_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_2_tile_v_6_1 = rf_matrix_b_2_tile_v_1_MPORT_6_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_2_tile_v_6_0 = rf_matrix_b_2_tile_v_0_MPORT_6_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_b_2_T_6 = {matrix_b_2_tile_v_6_3,matrix_b_2_tile_v_6_2,matrix_b_2_tile_v_6_1,
    matrix_b_2_tile_v_6_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] matrix_c_2_tile_v_6_3 = rf_matrix_c_2_tile_v_3_MPORT_6_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_2_tile_v_6_2 = rf_matrix_c_2_tile_v_2_MPORT_6_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_2_tile_v_6_1 = rf_matrix_c_2_tile_v_1_MPORT_6_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_2_tile_v_6_0 = rf_matrix_c_2_tile_v_0_MPORT_6_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_c_2_T_6 = {matrix_c_2_tile_v_6_3,matrix_c_2_tile_v_6_2,matrix_c_2_tile_v_6_1,
    matrix_c_2_tile_v_6_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] a_tile_v_55_3 = rf_a_tile_v_3_MPORT_18_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] a_tile_v_55_2 = rf_a_tile_v_2_MPORT_18_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] a_tile_v_55_1 = rf_a_tile_v_1_MPORT_55_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] a_tile_v_55_0 = rf_a_tile_v_0_MPORT_55_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] a_55 = {a_tile_v_55_3,a_tile_v_55_2,a_tile_v_55_1,a_tile_v_55_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] matrix_b_2_tile_v_7_3 = rf_matrix_b_2_tile_v_3_MPORT_7_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_2_tile_v_7_2 = rf_matrix_b_2_tile_v_2_MPORT_7_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_2_tile_v_7_1 = rf_matrix_b_2_tile_v_1_MPORT_7_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_2_tile_v_7_0 = rf_matrix_b_2_tile_v_0_MPORT_7_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_b_2_T_7 = {matrix_b_2_tile_v_7_3,matrix_b_2_tile_v_7_2,matrix_b_2_tile_v_7_1,
    matrix_b_2_tile_v_7_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] matrix_c_2_tile_v_7_3 = rf_matrix_c_2_tile_v_3_MPORT_7_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_2_tile_v_7_2 = rf_matrix_c_2_tile_v_2_MPORT_7_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_2_tile_v_7_1 = rf_matrix_c_2_tile_v_1_MPORT_7_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_2_tile_v_7_0 = rf_matrix_c_2_tile_v_0_MPORT_7_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_c_2_T_7 = {matrix_c_2_tile_v_7_3,matrix_c_2_tile_v_7_2,matrix_c_2_tile_v_7_1,
    matrix_c_2_tile_v_7_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [255:0] _GEN_3325 = io_mixPc ? _matrix_a_2_T_4 : a_55; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 256:30 258:29 263:29]
  wire [255:0] _GEN_3330 = io_mixPc ? _matrix_b_2_T_6 : _matrix_b_2_T_7; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 256:30 259:29 264:29]
  wire [255:0] _GEN_3331 = io_mixPc ? _matrix_c_2_T_6 : _matrix_c_2_T_7; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 256:30 260:29 265:29]
  wire [63:0] a_tile_v_56_1 = rf_a_tile_v_1_MPORT_56_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] a_tile_v_56_0 = rf_a_tile_v_0_MPORT_56_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_a_2_T_5 = {a_tile_v_56_1,a_tile_v_56_0,128'h0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 271:35]
  wire [63:0] matrix_b_2_tile_v_8_3 = rf_matrix_b_2_tile_v_3_MPORT_8_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_2_tile_v_8_2 = rf_matrix_b_2_tile_v_2_MPORT_8_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_2_tile_v_8_1 = rf_matrix_b_2_tile_v_1_MPORT_8_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_2_tile_v_8_0 = rf_matrix_b_2_tile_v_0_MPORT_8_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_b_2_T_8 = {matrix_b_2_tile_v_8_3,matrix_b_2_tile_v_8_2,matrix_b_2_tile_v_8_1,
    matrix_b_2_tile_v_8_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] matrix_c_2_tile_v_8_3 = rf_matrix_c_2_tile_v_3_MPORT_8_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_2_tile_v_8_2 = rf_matrix_c_2_tile_v_2_MPORT_8_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_2_tile_v_8_1 = rf_matrix_c_2_tile_v_1_MPORT_8_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_2_tile_v_8_0 = rf_matrix_c_2_tile_v_0_MPORT_8_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_c_2_T_8 = {matrix_c_2_tile_v_8_3,matrix_c_2_tile_v_8_2,matrix_c_2_tile_v_8_1,
    matrix_c_2_tile_v_8_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] a_tile_v_57_3 = rf_a_tile_v_3_MPORT_19_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] a_tile_v_57_2 = rf_a_tile_v_2_MPORT_19_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] a_tile_v_57_1 = rf_a_tile_v_1_MPORT_57_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] a_tile_v_57_0 = rf_a_tile_v_0_MPORT_57_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] a_57 = {a_tile_v_57_3,a_tile_v_57_2,a_tile_v_57_1,a_tile_v_57_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] matrix_b_2_tile_v_9_3 = rf_matrix_b_2_tile_v_3_MPORT_9_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_2_tile_v_9_2 = rf_matrix_b_2_tile_v_2_MPORT_9_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_2_tile_v_9_1 = rf_matrix_b_2_tile_v_1_MPORT_9_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_2_tile_v_9_0 = rf_matrix_b_2_tile_v_0_MPORT_9_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_b_2_T_9 = {matrix_b_2_tile_v_9_3,matrix_b_2_tile_v_9_2,matrix_b_2_tile_v_9_1,
    matrix_b_2_tile_v_9_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] matrix_c_2_tile_v_9_3 = rf_matrix_c_2_tile_v_3_MPORT_9_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_2_tile_v_9_2 = rf_matrix_c_2_tile_v_2_MPORT_9_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_2_tile_v_9_1 = rf_matrix_c_2_tile_v_1_MPORT_9_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_2_tile_v_9_0 = rf_matrix_c_2_tile_v_0_MPORT_9_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_c_2_T_9 = {matrix_c_2_tile_v_9_3,matrix_c_2_tile_v_9_2,matrix_c_2_tile_v_9_1,
    matrix_c_2_tile_v_9_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [255:0] _GEN_3336 = io_mixPc ? _matrix_a_2_T_5 : a_57; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 269:30 271:29 276:29]
  wire [255:0] _GEN_3337 = io_mixPc ? _matrix_b_2_T_8 : _matrix_b_2_T_9; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 269:30 272:29 277:29]
  wire [255:0] _GEN_3338 = io_mixPc ? _matrix_c_2_T_8 : _matrix_c_2_T_9; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 269:30 273:29 278:29]
  wire [63:0] a_tile_v_58_1 = rf_a_tile_v_1_MPORT_58_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] a_tile_v_58_0 = rf_a_tile_v_0_MPORT_58_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_a_2_T_6 = {a_tile_v_58_1,a_tile_v_58_0,128'h0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 283:33]
  wire [63:0] matrix_b_2_tile_v_10_3 = rf_matrix_b_2_tile_v_3_MPORT_10_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_2_tile_v_10_2 = rf_matrix_b_2_tile_v_2_MPORT_10_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_2_tile_v_10_1 = rf_matrix_b_2_tile_v_1_MPORT_10_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_2_tile_v_10_0 = rf_matrix_b_2_tile_v_0_MPORT_10_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_b_2_T_10 = {matrix_b_2_tile_v_10_3,matrix_b_2_tile_v_10_2,matrix_b_2_tile_v_10_1,
    matrix_b_2_tile_v_10_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] matrix_c_2_tile_v_10_3 = rf_matrix_c_2_tile_v_3_MPORT_10_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_2_tile_v_10_2 = rf_matrix_c_2_tile_v_2_MPORT_10_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_2_tile_v_10_1 = rf_matrix_c_2_tile_v_1_MPORT_10_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_2_tile_v_10_0 = rf_matrix_c_2_tile_v_0_MPORT_10_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_c_2_T_10 = {matrix_c_2_tile_v_10_3,matrix_c_2_tile_v_10_2,matrix_c_2_tile_v_10_1,
    matrix_c_2_tile_v_10_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] a_tile_v_59_1 = rf_a_tile_v_1_MPORT_59_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] a_tile_v_59_0 = rf_a_tile_v_0_MPORT_59_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_a_2_T_7 = {a_tile_v_59_1,a_tile_v_59_0,128'h0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 289:33]
  wire [63:0] matrix_b_2_tile_v_11_3 = rf_matrix_b_2_tile_v_3_MPORT_11_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_2_tile_v_11_2 = rf_matrix_b_2_tile_v_2_MPORT_11_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_2_tile_v_11_1 = rf_matrix_b_2_tile_v_1_MPORT_11_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_2_tile_v_11_0 = rf_matrix_b_2_tile_v_0_MPORT_11_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_b_2_T_11 = {matrix_b_2_tile_v_11_3,matrix_b_2_tile_v_11_2,matrix_b_2_tile_v_11_1,
    matrix_b_2_tile_v_11_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] matrix_c_2_tile_v_11_3 = rf_matrix_c_2_tile_v_3_MPORT_11_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_2_tile_v_11_2 = rf_matrix_c_2_tile_v_2_MPORT_11_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_2_tile_v_11_1 = rf_matrix_c_2_tile_v_1_MPORT_11_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_2_tile_v_11_0 = rf_matrix_c_2_tile_v_0_MPORT_11_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_c_2_T_11 = {matrix_c_2_tile_v_11_3,matrix_c_2_tile_v_11_2,matrix_c_2_tile_v_11_1,
    matrix_c_2_tile_v_11_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [255:0] _GEN_3343 = _T_4 ? _matrix_a_2_T_7 : matrix_a_2; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 159:21 254:24 289:27]
  wire [255:0] _GEN_3348 = _T_4 ? _matrix_b_2_T_11 : matrix_b_2; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 160:21 254:24 290:27]
  wire [255:0] _GEN_3353 = _T_4 ? _matrix_c_2_T_11 : matrix_c_2; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 161:21 254:24 291:27]
  wire [255:0] _GEN_3358 = _T_3 ? _matrix_a_2_T_6 : _GEN_3343; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 254:24 283:27]
  wire [255:0] _GEN_3363 = _T_3 ? _matrix_b_2_T_10 : _GEN_3348; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 254:24 284:27]
  wire [255:0] _GEN_3368 = _T_3 ? _matrix_c_2_T_10 : _GEN_3353; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 254:24 285:27]
  wire [255:0] _GEN_3385 = _T_2 ? _GEN_3336 : _GEN_3358; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 254:24]
  wire [255:0] _GEN_3390 = _T_2 ? _GEN_3337 : _GEN_3363; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 254:24]
  wire [255:0] _GEN_3395 = _T_2 ? _GEN_3338 : _GEN_3368; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 254:24]
  wire [63:0] a_tile_v_60_1 = rf_a_tile_v_1_MPORT_60_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] a_tile_v_60_0 = rf_a_tile_v_0_MPORT_60_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_a_2_T_8 = {a_tile_v_60_1,a_tile_v_60_0,128'h0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 300:35]
  wire [63:0] matrix_b_2_tile_v_12_3 = rf_matrix_b_2_tile_v_3_MPORT_12_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_2_tile_v_12_2 = rf_matrix_b_2_tile_v_2_MPORT_12_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_2_tile_v_12_1 = rf_matrix_b_2_tile_v_1_MPORT_12_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_2_tile_v_12_0 = rf_matrix_b_2_tile_v_0_MPORT_12_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_b_2_T_12 = {matrix_b_2_tile_v_12_3,matrix_b_2_tile_v_12_2,matrix_b_2_tile_v_12_1,
    matrix_b_2_tile_v_12_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] matrix_c_2_tile_v_12_3 = rf_matrix_c_2_tile_v_3_MPORT_12_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_2_tile_v_12_2 = rf_matrix_c_2_tile_v_2_MPORT_12_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_2_tile_v_12_1 = rf_matrix_c_2_tile_v_1_MPORT_12_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_2_tile_v_12_0 = rf_matrix_c_2_tile_v_0_MPORT_12_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_c_2_T_12 = {matrix_c_2_tile_v_12_3,matrix_c_2_tile_v_12_2,matrix_c_2_tile_v_12_1,
    matrix_c_2_tile_v_12_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] a_tile_v_61_3 = rf_a_tile_v_3_MPORT_20_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] a_tile_v_61_2 = rf_a_tile_v_2_MPORT_20_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] a_tile_v_61_1 = rf_a_tile_v_1_MPORT_61_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] a_tile_v_61_0 = rf_a_tile_v_0_MPORT_61_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] a_61 = {a_tile_v_61_3,a_tile_v_61_2,a_tile_v_61_1,a_tile_v_61_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] matrix_b_2_tile_v_13_3 = rf_matrix_b_2_tile_v_3_MPORT_13_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_2_tile_v_13_2 = rf_matrix_b_2_tile_v_2_MPORT_13_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_2_tile_v_13_1 = rf_matrix_b_2_tile_v_1_MPORT_13_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_2_tile_v_13_0 = rf_matrix_b_2_tile_v_0_MPORT_13_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_b_2_T_13 = {matrix_b_2_tile_v_13_3,matrix_b_2_tile_v_13_2,matrix_b_2_tile_v_13_1,
    matrix_b_2_tile_v_13_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] matrix_c_2_tile_v_13_3 = rf_matrix_c_2_tile_v_3_MPORT_13_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_2_tile_v_13_2 = rf_matrix_c_2_tile_v_2_MPORT_13_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_2_tile_v_13_1 = rf_matrix_c_2_tile_v_1_MPORT_13_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_2_tile_v_13_0 = rf_matrix_c_2_tile_v_0_MPORT_13_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_c_2_T_13 = {matrix_c_2_tile_v_13_3,matrix_c_2_tile_v_13_2,matrix_c_2_tile_v_13_1,
    matrix_c_2_tile_v_13_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [255:0] _GEN_3513 = io_mixPc ? _matrix_a_2_T_8 : a_61; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 298:30 300:29 305:29]
  wire [255:0] _GEN_3518 = io_mixPc ? _matrix_b_2_T_12 : _matrix_b_2_T_13; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 298:30 301:29 306:29]
  wire [255:0] _GEN_3519 = io_mixPc ? _matrix_c_2_T_12 : _matrix_c_2_T_13; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 298:30 302:29 307:29]
  wire [63:0] a_tile_v_62_1 = rf_a_tile_v_1_MPORT_62_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] a_tile_v_62_0 = rf_a_tile_v_0_MPORT_62_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_a_2_T_9 = {a_tile_v_62_1,a_tile_v_62_0,128'h0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 313:35]
  wire [63:0] matrix_b_2_tile_v_14_3 = rf_matrix_b_2_tile_v_3_MPORT_14_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_2_tile_v_14_2 = rf_matrix_b_2_tile_v_2_MPORT_14_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_2_tile_v_14_1 = rf_matrix_b_2_tile_v_1_MPORT_14_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_2_tile_v_14_0 = rf_matrix_b_2_tile_v_0_MPORT_14_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_b_2_T_14 = {matrix_b_2_tile_v_14_3,matrix_b_2_tile_v_14_2,matrix_b_2_tile_v_14_1,
    matrix_b_2_tile_v_14_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] matrix_c_2_tile_v_14_3 = rf_matrix_c_2_tile_v_3_MPORT_14_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_2_tile_v_14_2 = rf_matrix_c_2_tile_v_2_MPORT_14_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_2_tile_v_14_1 = rf_matrix_c_2_tile_v_1_MPORT_14_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_2_tile_v_14_0 = rf_matrix_c_2_tile_v_0_MPORT_14_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_c_2_T_14 = {matrix_c_2_tile_v_14_3,matrix_c_2_tile_v_14_2,matrix_c_2_tile_v_14_1,
    matrix_c_2_tile_v_14_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] a_tile_v_63_3 = rf_a_tile_v_3_MPORT_21_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] a_tile_v_63_2 = rf_a_tile_v_2_MPORT_21_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] a_tile_v_63_1 = rf_a_tile_v_1_MPORT_63_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] a_tile_v_63_0 = rf_a_tile_v_0_MPORT_63_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] a_63 = {a_tile_v_63_3,a_tile_v_63_2,a_tile_v_63_1,a_tile_v_63_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] matrix_b_2_tile_v_15_3 = rf_matrix_b_2_tile_v_3_MPORT_15_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_2_tile_v_15_2 = rf_matrix_b_2_tile_v_2_MPORT_15_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_2_tile_v_15_1 = rf_matrix_b_2_tile_v_1_MPORT_15_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_2_tile_v_15_0 = rf_matrix_b_2_tile_v_0_MPORT_15_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_b_2_T_15 = {matrix_b_2_tile_v_15_3,matrix_b_2_tile_v_15_2,matrix_b_2_tile_v_15_1,
    matrix_b_2_tile_v_15_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] matrix_c_2_tile_v_15_3 = rf_matrix_c_2_tile_v_3_MPORT_15_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_2_tile_v_15_2 = rf_matrix_c_2_tile_v_2_MPORT_15_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_2_tile_v_15_1 = rf_matrix_c_2_tile_v_1_MPORT_15_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_2_tile_v_15_0 = rf_matrix_c_2_tile_v_0_MPORT_15_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_c_2_T_15 = {matrix_c_2_tile_v_15_3,matrix_c_2_tile_v_15_2,matrix_c_2_tile_v_15_1,
    matrix_c_2_tile_v_15_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [255:0] _GEN_3524 = io_mixPc ? _matrix_a_2_T_9 : a_63; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 311:30 313:29 318:29]
  wire [255:0] _GEN_3525 = io_mixPc ? _matrix_b_2_T_14 : _matrix_b_2_T_15; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 311:30 314:29 319:29]
  wire [255:0] _GEN_3526 = io_mixPc ? _matrix_c_2_T_14 : _matrix_c_2_T_15; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 311:30 315:29 320:29]
  wire [63:0] a_tile_v_64_1 = rf_a_tile_v_1_MPORT_64_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] a_tile_v_64_0 = rf_a_tile_v_0_MPORT_64_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_a_2_T_10 = {a_tile_v_64_1,a_tile_v_64_0,128'h0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 325:33]
  wire [63:0] matrix_b_2_tile_v_16_3 = rf_matrix_b_2_tile_v_3_MPORT_16_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_2_tile_v_16_2 = rf_matrix_b_2_tile_v_2_MPORT_16_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_2_tile_v_16_1 = rf_matrix_b_2_tile_v_1_MPORT_16_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_2_tile_v_16_0 = rf_matrix_b_2_tile_v_0_MPORT_16_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_b_2_T_16 = {matrix_b_2_tile_v_16_3,matrix_b_2_tile_v_16_2,matrix_b_2_tile_v_16_1,
    matrix_b_2_tile_v_16_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] matrix_c_2_tile_v_16_3 = rf_matrix_c_2_tile_v_3_MPORT_16_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_2_tile_v_16_2 = rf_matrix_c_2_tile_v_2_MPORT_16_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_2_tile_v_16_1 = rf_matrix_c_2_tile_v_1_MPORT_16_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_2_tile_v_16_0 = rf_matrix_c_2_tile_v_0_MPORT_16_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_c_2_T_16 = {matrix_c_2_tile_v_16_3,matrix_c_2_tile_v_16_2,matrix_c_2_tile_v_16_1,
    matrix_c_2_tile_v_16_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] a_tile_v_65_1 = rf_a_tile_v_1_MPORT_65_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] a_tile_v_65_0 = rf_a_tile_v_0_MPORT_65_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_a_2_T_11 = {a_tile_v_65_1,a_tile_v_65_0,128'h0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 331:33]
  wire [63:0] matrix_b_2_tile_v_17_3 = rf_matrix_b_2_tile_v_3_MPORT_17_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_2_tile_v_17_2 = rf_matrix_b_2_tile_v_2_MPORT_17_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_2_tile_v_17_1 = rf_matrix_b_2_tile_v_1_MPORT_17_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_2_tile_v_17_0 = rf_matrix_b_2_tile_v_0_MPORT_17_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_b_2_T_17 = {matrix_b_2_tile_v_17_3,matrix_b_2_tile_v_17_2,matrix_b_2_tile_v_17_1,
    matrix_b_2_tile_v_17_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] matrix_c_2_tile_v_17_3 = rf_matrix_c_2_tile_v_3_MPORT_17_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_2_tile_v_17_2 = rf_matrix_c_2_tile_v_2_MPORT_17_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_2_tile_v_17_1 = rf_matrix_c_2_tile_v_1_MPORT_17_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_2_tile_v_17_0 = rf_matrix_c_2_tile_v_0_MPORT_17_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_c_2_T_17 = {matrix_c_2_tile_v_17_3,matrix_c_2_tile_v_17_2,matrix_c_2_tile_v_17_1,
    matrix_c_2_tile_v_17_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [255:0] _GEN_3531 = _T_4 ? _matrix_a_2_T_11 : matrix_a_2; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 159:21 296:24 331:27]
  wire [255:0] _GEN_3536 = _T_4 ? _matrix_b_2_T_17 : matrix_b_2; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 160:21 296:24 332:27]
  wire [255:0] _GEN_3541 = _T_4 ? _matrix_c_2_T_17 : matrix_c_2; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 161:21 296:24 333:27]
  wire [255:0] _GEN_3546 = _T_3 ? _matrix_a_2_T_10 : _GEN_3531; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 296:24 325:27]
  wire [255:0] _GEN_3551 = _T_3 ? _matrix_b_2_T_16 : _GEN_3536; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 296:24 326:27]
  wire [255:0] _GEN_3556 = _T_3 ? _matrix_c_2_T_16 : _GEN_3541; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 296:24 327:27]
  wire [255:0] _GEN_3573 = _T_2 ? _GEN_3524 : _GEN_3546; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 296:24]
  wire [255:0] _GEN_3578 = _T_2 ? _GEN_3525 : _GEN_3551; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 296:24]
  wire [255:0] _GEN_3583 = _T_2 ? _GEN_3526 : _GEN_3556; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 296:24]
  wire [255:0] _GEN_3626 = _T_1 ? _GEN_3513 : _GEN_3573; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 296:24]
  wire [255:0] _GEN_3631 = _T_1 ? _GEN_3518 : _GEN_3578; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 296:24]
  wire [255:0] _GEN_3636 = _T_1 ? _GEN_3519 : _GEN_3583; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 296:24]
  wire [63:0] a_tile_v_66_1 = rf_a_tile_v_1_MPORT_66_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] a_tile_v_66_0 = rf_a_tile_v_0_MPORT_66_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_a_2_T_12 = {a_tile_v_66_1,a_tile_v_66_0,128'h0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 342:35]
  wire [63:0] matrix_b_2_tile_v_18_3 = rf_matrix_b_2_tile_v_3_MPORT_18_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_2_tile_v_18_2 = rf_matrix_b_2_tile_v_2_MPORT_18_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_2_tile_v_18_1 = rf_matrix_b_2_tile_v_1_MPORT_18_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_2_tile_v_18_0 = rf_matrix_b_2_tile_v_0_MPORT_18_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_b_2_T_18 = {matrix_b_2_tile_v_18_3,matrix_b_2_tile_v_18_2,matrix_b_2_tile_v_18_1,
    matrix_b_2_tile_v_18_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] matrix_c_2_tile_v_18_3 = rf_matrix_c_2_tile_v_3_MPORT_18_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_2_tile_v_18_2 = rf_matrix_c_2_tile_v_2_MPORT_18_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_2_tile_v_18_1 = rf_matrix_c_2_tile_v_1_MPORT_18_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_2_tile_v_18_0 = rf_matrix_c_2_tile_v_0_MPORT_18_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_c_2_T_18 = {matrix_c_2_tile_v_18_3,matrix_c_2_tile_v_18_2,matrix_c_2_tile_v_18_1,
    matrix_c_2_tile_v_18_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] a_tile_v_67_3 = rf_a_tile_v_3_MPORT_22_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] a_tile_v_67_2 = rf_a_tile_v_2_MPORT_22_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] a_tile_v_67_1 = rf_a_tile_v_1_MPORT_67_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] a_tile_v_67_0 = rf_a_tile_v_0_MPORT_67_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] a_67 = {a_tile_v_67_3,a_tile_v_67_2,a_tile_v_67_1,a_tile_v_67_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] matrix_b_2_tile_v_19_3 = rf_matrix_b_2_tile_v_3_MPORT_19_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_2_tile_v_19_2 = rf_matrix_b_2_tile_v_2_MPORT_19_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_2_tile_v_19_1 = rf_matrix_b_2_tile_v_1_MPORT_19_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_2_tile_v_19_0 = rf_matrix_b_2_tile_v_0_MPORT_19_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_b_2_T_19 = {matrix_b_2_tile_v_19_3,matrix_b_2_tile_v_19_2,matrix_b_2_tile_v_19_1,
    matrix_b_2_tile_v_19_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] matrix_c_2_tile_v_19_3 = rf_matrix_c_2_tile_v_3_MPORT_19_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_2_tile_v_19_2 = rf_matrix_c_2_tile_v_2_MPORT_19_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_2_tile_v_19_1 = rf_matrix_c_2_tile_v_1_MPORT_19_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_2_tile_v_19_0 = rf_matrix_c_2_tile_v_0_MPORT_19_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_c_2_T_19 = {matrix_c_2_tile_v_19_3,matrix_c_2_tile_v_19_2,matrix_c_2_tile_v_19_1,
    matrix_c_2_tile_v_19_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [255:0] _GEN_3701 = io_mixPc ? _matrix_a_2_T_12 : a_67; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 340:30 342:29 347:29]
  wire [255:0] _GEN_3706 = io_mixPc ? _matrix_b_2_T_18 : _matrix_b_2_T_19; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 340:30 343:29 348:29]
  wire [255:0] _GEN_3707 = io_mixPc ? _matrix_c_2_T_18 : _matrix_c_2_T_19; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 340:30 344:29 349:29]
  wire [63:0] a_tile_v_68_1 = rf_a_tile_v_1_MPORT_68_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] a_tile_v_68_0 = rf_a_tile_v_0_MPORT_68_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_a_2_T_13 = {a_tile_v_68_1,a_tile_v_68_0,128'h0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 355:35]
  wire [63:0] matrix_b_2_tile_v_20_3 = rf_matrix_b_2_tile_v_3_MPORT_20_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_2_tile_v_20_2 = rf_matrix_b_2_tile_v_2_MPORT_20_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_2_tile_v_20_1 = rf_matrix_b_2_tile_v_1_MPORT_20_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_2_tile_v_20_0 = rf_matrix_b_2_tile_v_0_MPORT_20_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_b_2_T_20 = {matrix_b_2_tile_v_20_3,matrix_b_2_tile_v_20_2,matrix_b_2_tile_v_20_1,
    matrix_b_2_tile_v_20_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] matrix_c_2_tile_v_20_3 = rf_matrix_c_2_tile_v_3_MPORT_20_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_2_tile_v_20_2 = rf_matrix_c_2_tile_v_2_MPORT_20_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_2_tile_v_20_1 = rf_matrix_c_2_tile_v_1_MPORT_20_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_2_tile_v_20_0 = rf_matrix_c_2_tile_v_0_MPORT_20_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_c_2_T_20 = {matrix_c_2_tile_v_20_3,matrix_c_2_tile_v_20_2,matrix_c_2_tile_v_20_1,
    matrix_c_2_tile_v_20_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] a_tile_v_69_3 = rf_a_tile_v_3_MPORT_23_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] a_tile_v_69_2 = rf_a_tile_v_2_MPORT_23_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] a_tile_v_69_1 = rf_a_tile_v_1_MPORT_69_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] a_tile_v_69_0 = rf_a_tile_v_0_MPORT_69_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] a_69 = {a_tile_v_69_3,a_tile_v_69_2,a_tile_v_69_1,a_tile_v_69_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] matrix_b_2_tile_v_21_3 = rf_matrix_b_2_tile_v_3_MPORT_21_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_2_tile_v_21_2 = rf_matrix_b_2_tile_v_2_MPORT_21_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_2_tile_v_21_1 = rf_matrix_b_2_tile_v_1_MPORT_21_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_2_tile_v_21_0 = rf_matrix_b_2_tile_v_0_MPORT_21_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_b_2_T_21 = {matrix_b_2_tile_v_21_3,matrix_b_2_tile_v_21_2,matrix_b_2_tile_v_21_1,
    matrix_b_2_tile_v_21_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] matrix_c_2_tile_v_21_3 = rf_matrix_c_2_tile_v_3_MPORT_21_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_2_tile_v_21_2 = rf_matrix_c_2_tile_v_2_MPORT_21_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_2_tile_v_21_1 = rf_matrix_c_2_tile_v_1_MPORT_21_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_2_tile_v_21_0 = rf_matrix_c_2_tile_v_0_MPORT_21_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_c_2_T_21 = {matrix_c_2_tile_v_21_3,matrix_c_2_tile_v_21_2,matrix_c_2_tile_v_21_1,
    matrix_c_2_tile_v_21_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [255:0] _GEN_3712 = io_mixPc ? _matrix_a_2_T_13 : a_69; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 353:30 355:29 360:29]
  wire [255:0] _GEN_3713 = io_mixPc ? _matrix_b_2_T_20 : _matrix_b_2_T_21; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 353:30 356:29 361:29]
  wire [255:0] _GEN_3714 = io_mixPc ? _matrix_c_2_T_20 : _matrix_c_2_T_21; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 353:30 357:29 362:29]
  wire [63:0] a_tile_v_70_1 = rf_a_tile_v_1_MPORT_70_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] a_tile_v_70_0 = rf_a_tile_v_0_MPORT_70_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_a_2_T_14 = {a_tile_v_70_1,a_tile_v_70_0,128'h0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 367:33]
  wire [63:0] matrix_b_2_tile_v_22_3 = rf_matrix_b_2_tile_v_3_MPORT_22_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_2_tile_v_22_2 = rf_matrix_b_2_tile_v_2_MPORT_22_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_2_tile_v_22_1 = rf_matrix_b_2_tile_v_1_MPORT_22_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_2_tile_v_22_0 = rf_matrix_b_2_tile_v_0_MPORT_22_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_b_2_T_22 = {matrix_b_2_tile_v_22_3,matrix_b_2_tile_v_22_2,matrix_b_2_tile_v_22_1,
    matrix_b_2_tile_v_22_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] matrix_c_2_tile_v_22_3 = rf_matrix_c_2_tile_v_3_MPORT_22_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_2_tile_v_22_2 = rf_matrix_c_2_tile_v_2_MPORT_22_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_2_tile_v_22_1 = rf_matrix_c_2_tile_v_1_MPORT_22_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_2_tile_v_22_0 = rf_matrix_c_2_tile_v_0_MPORT_22_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_c_2_T_22 = {matrix_c_2_tile_v_22_3,matrix_c_2_tile_v_22_2,matrix_c_2_tile_v_22_1,
    matrix_c_2_tile_v_22_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] a_tile_v_71_1 = rf_a_tile_v_1_MPORT_71_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] a_tile_v_71_0 = rf_a_tile_v_0_MPORT_71_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_a_2_T_15 = {a_tile_v_71_1,a_tile_v_71_0,128'h0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 373:33]
  wire [63:0] matrix_b_2_tile_v_23_3 = rf_matrix_b_2_tile_v_3_MPORT_23_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_2_tile_v_23_2 = rf_matrix_b_2_tile_v_2_MPORT_23_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_2_tile_v_23_1 = rf_matrix_b_2_tile_v_1_MPORT_23_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_2_tile_v_23_0 = rf_matrix_b_2_tile_v_0_MPORT_23_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_b_2_T_23 = {matrix_b_2_tile_v_23_3,matrix_b_2_tile_v_23_2,matrix_b_2_tile_v_23_1,
    matrix_b_2_tile_v_23_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] matrix_c_2_tile_v_23_3 = rf_matrix_c_2_tile_v_3_MPORT_23_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_2_tile_v_23_2 = rf_matrix_c_2_tile_v_2_MPORT_23_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_2_tile_v_23_1 = rf_matrix_c_2_tile_v_1_MPORT_23_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_2_tile_v_23_0 = rf_matrix_c_2_tile_v_0_MPORT_23_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_c_2_T_23 = {matrix_c_2_tile_v_23_3,matrix_c_2_tile_v_23_2,matrix_c_2_tile_v_23_1,
    matrix_c_2_tile_v_23_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [255:0] _GEN_3719 = _T_4 ? _matrix_a_2_T_15 : matrix_a_2; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 159:21 338:24 373:27]
  wire [255:0] _GEN_3724 = _T_4 ? _matrix_b_2_T_23 : matrix_b_2; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 160:21 338:24 374:27]
  wire [255:0] _GEN_3729 = _T_4 ? _matrix_c_2_T_23 : matrix_c_2; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 161:21 338:24 375:27]
  wire [255:0] _GEN_3734 = _T_3 ? _matrix_a_2_T_14 : _GEN_3719; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 338:24 367:27]
  wire [255:0] _GEN_3739 = _T_3 ? _matrix_b_2_T_22 : _GEN_3724; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 338:24 368:27]
  wire [255:0] _GEN_3744 = _T_3 ? _matrix_c_2_T_22 : _GEN_3729; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 338:24 369:27]
  wire [255:0] _GEN_3761 = _T_2 ? _GEN_3712 : _GEN_3734; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 338:24]
  wire [255:0] _GEN_3766 = _T_2 ? _GEN_3713 : _GEN_3739; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 338:24]
  wire [255:0] _GEN_3771 = _T_2 ? _GEN_3714 : _GEN_3744; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 338:24]
  wire [255:0] _GEN_3814 = _T_1 ? _GEN_3701 : _GEN_3761; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 338:24]
  wire [255:0] _GEN_3819 = _T_1 ? _GEN_3706 : _GEN_3766; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 338:24]
  wire [255:0] _GEN_3824 = _T_1 ? _GEN_3707 : _GEN_3771; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 338:24]
  wire [255:0] _GEN_3893 = 2'h3 == set ? _GEN_3814 : matrix_a_2; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 210:18 159:21]
  wire [255:0] _GEN_3898 = 2'h3 == set ? _GEN_3819 : matrix_b_2; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 210:18 160:21]
  wire [255:0] _GEN_3903 = 2'h3 == set ? _GEN_3824 : matrix_c_2; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 210:18 161:21]
  wire [63:0] a_tile_v_72_1 = rf_a_tile_v_1_MPORT_72_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] a_tile_v_72_0 = rf_a_tile_v_0_MPORT_72_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_a_3_T = {a_tile_v_72_1,a_tile_v_72_0,128'h0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 216:35]
  wire [63:0] matrix_b_3_tile_v__3 = rf_matrix_b_3_tile_v_3_MPORT_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_3_tile_v__2 = rf_matrix_b_3_tile_v_2_MPORT_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_3_tile_v__1 = rf_matrix_b_3_tile_v_1_MPORT_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_3_tile_v__0 = rf_matrix_b_3_tile_v_0_MPORT_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_b_3_T = {matrix_b_3_tile_v__3,matrix_b_3_tile_v__2,matrix_b_3_tile_v__1,matrix_b_3_tile_v__0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] matrix_c_3_tile_v__3 = rf_matrix_c_3_tile_v_3_MPORT_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_3_tile_v__2 = rf_matrix_c_3_tile_v_2_MPORT_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_3_tile_v__1 = rf_matrix_c_3_tile_v_1_MPORT_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_3_tile_v__0 = rf_matrix_c_3_tile_v_0_MPORT_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_c_3_T = {matrix_c_3_tile_v__3,matrix_c_3_tile_v__2,matrix_c_3_tile_v__1,matrix_c_3_tile_v__0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] a_tile_v_73_3 = rf_a_tile_v_3_MPORT_24_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] a_tile_v_73_2 = rf_a_tile_v_2_MPORT_24_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] a_tile_v_73_1 = rf_a_tile_v_1_MPORT_73_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] a_tile_v_73_0 = rf_a_tile_v_0_MPORT_73_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] a_73 = {a_tile_v_73_3,a_tile_v_73_2,a_tile_v_73_1,a_tile_v_73_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] matrix_b_3_tile_v_1_3 = rf_matrix_b_3_tile_v_3_MPORT_1_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_3_tile_v_1_2 = rf_matrix_b_3_tile_v_2_MPORT_1_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_3_tile_v_1_1 = rf_matrix_b_3_tile_v_1_MPORT_1_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_3_tile_v_1_0 = rf_matrix_b_3_tile_v_0_MPORT_1_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_b_3_T_1 = {matrix_b_3_tile_v_1_3,matrix_b_3_tile_v_1_2,matrix_b_3_tile_v_1_1,
    matrix_b_3_tile_v_1_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] matrix_c_3_tile_v_1_3 = rf_matrix_c_3_tile_v_3_MPORT_1_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_3_tile_v_1_2 = rf_matrix_c_3_tile_v_2_MPORT_1_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_3_tile_v_1_1 = rf_matrix_c_3_tile_v_1_MPORT_1_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_3_tile_v_1_0 = rf_matrix_c_3_tile_v_0_MPORT_1_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_c_3_T_1 = {matrix_c_3_tile_v_1_3,matrix_c_3_tile_v_1_2,matrix_c_3_tile_v_1_1,
    matrix_c_3_tile_v_1_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] a_tile_v_74_1 = rf_a_tile_v_1_MPORT_74_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] a_tile_v_74_0 = rf_a_tile_v_0_MPORT_74_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_a_3_T_1 = {a_tile_v_74_1,a_tile_v_74_0,128'h0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 229:35]
  wire [63:0] matrix_b_3_tile_v_2_3 = rf_matrix_b_3_tile_v_3_MPORT_2_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_3_tile_v_2_2 = rf_matrix_b_3_tile_v_2_MPORT_2_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_3_tile_v_2_1 = rf_matrix_b_3_tile_v_1_MPORT_2_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_3_tile_v_2_0 = rf_matrix_b_3_tile_v_0_MPORT_2_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_b_3_T_2 = {matrix_b_3_tile_v_2_3,matrix_b_3_tile_v_2_2,matrix_b_3_tile_v_2_1,
    matrix_b_3_tile_v_2_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] matrix_c_3_tile_v_2_3 = rf_matrix_c_3_tile_v_3_MPORT_2_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_3_tile_v_2_2 = rf_matrix_c_3_tile_v_2_MPORT_2_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_3_tile_v_2_1 = rf_matrix_c_3_tile_v_1_MPORT_2_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_3_tile_v_2_0 = rf_matrix_c_3_tile_v_0_MPORT_2_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_c_3_T_2 = {matrix_c_3_tile_v_2_3,matrix_c_3_tile_v_2_2,matrix_c_3_tile_v_2_1,
    matrix_c_3_tile_v_2_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] a_tile_v_75_3 = rf_a_tile_v_3_MPORT_25_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] a_tile_v_75_2 = rf_a_tile_v_2_MPORT_25_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] a_tile_v_75_1 = rf_a_tile_v_1_MPORT_75_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] a_tile_v_75_0 = rf_a_tile_v_0_MPORT_75_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] a_75 = {a_tile_v_75_3,a_tile_v_75_2,a_tile_v_75_1,a_tile_v_75_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] matrix_b_3_tile_v_3_3 = rf_matrix_b_3_tile_v_3_MPORT_3_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_3_tile_v_3_2 = rf_matrix_b_3_tile_v_2_MPORT_3_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_3_tile_v_3_1 = rf_matrix_b_3_tile_v_1_MPORT_3_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_3_tile_v_3_0 = rf_matrix_b_3_tile_v_0_MPORT_3_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_b_3_T_3 = {matrix_b_3_tile_v_3_3,matrix_b_3_tile_v_3_2,matrix_b_3_tile_v_3_1,
    matrix_b_3_tile_v_3_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] matrix_c_3_tile_v_3_3 = rf_matrix_c_3_tile_v_3_MPORT_3_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_3_tile_v_3_2 = rf_matrix_c_3_tile_v_2_MPORT_3_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_3_tile_v_3_1 = rf_matrix_c_3_tile_v_1_MPORT_3_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_3_tile_v_3_0 = rf_matrix_c_3_tile_v_0_MPORT_3_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_c_3_T_3 = {matrix_c_3_tile_v_3_3,matrix_c_3_tile_v_3_2,matrix_c_3_tile_v_3_1,
    matrix_c_3_tile_v_3_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [255:0] _GEN_4672 = io_mixPc ? _matrix_a_3_T_1 : a_75; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 227:30 229:29 234:29]
  wire [255:0] _GEN_4673 = io_mixPc ? _matrix_b_3_T_2 : _matrix_b_3_T_3; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 227:30 230:29 235:29]
  wire [255:0] _GEN_4678 = io_mixPc ? _matrix_c_3_T_2 : _matrix_c_3_T_3; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 227:30 231:29 236:29]
  wire [63:0] a_tile_v_76_1 = rf_a_tile_v_1_MPORT_76_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] a_tile_v_76_0 = rf_a_tile_v_0_MPORT_76_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_a_3_T_2 = {a_tile_v_76_1,a_tile_v_76_0,128'h0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 241:33]
  wire [63:0] matrix_b_3_tile_v_4_3 = rf_matrix_b_3_tile_v_3_MPORT_4_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_3_tile_v_4_2 = rf_matrix_b_3_tile_v_2_MPORT_4_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_3_tile_v_4_1 = rf_matrix_b_3_tile_v_1_MPORT_4_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_3_tile_v_4_0 = rf_matrix_b_3_tile_v_0_MPORT_4_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_b_3_T_4 = {matrix_b_3_tile_v_4_3,matrix_b_3_tile_v_4_2,matrix_b_3_tile_v_4_1,
    matrix_b_3_tile_v_4_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] matrix_c_3_tile_v_4_3 = rf_matrix_c_3_tile_v_3_MPORT_4_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_3_tile_v_4_2 = rf_matrix_c_3_tile_v_2_MPORT_4_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_3_tile_v_4_1 = rf_matrix_c_3_tile_v_1_MPORT_4_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_3_tile_v_4_0 = rf_matrix_c_3_tile_v_0_MPORT_4_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_c_3_T_4 = {matrix_c_3_tile_v_4_3,matrix_c_3_tile_v_4_2,matrix_c_3_tile_v_4_1,
    matrix_c_3_tile_v_4_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] a_tile_v_77_1 = rf_a_tile_v_1_MPORT_77_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] a_tile_v_77_0 = rf_a_tile_v_0_MPORT_77_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_a_3_T_3 = {a_tile_v_77_1,a_tile_v_77_0,128'h0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 247:33]
  wire [63:0] matrix_b_3_tile_v_5_3 = rf_matrix_b_3_tile_v_3_MPORT_5_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_3_tile_v_5_2 = rf_matrix_b_3_tile_v_2_MPORT_5_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_3_tile_v_5_1 = rf_matrix_b_3_tile_v_1_MPORT_5_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_3_tile_v_5_0 = rf_matrix_b_3_tile_v_0_MPORT_5_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_b_3_T_5 = {matrix_b_3_tile_v_5_3,matrix_b_3_tile_v_5_2,matrix_b_3_tile_v_5_1,
    matrix_b_3_tile_v_5_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] matrix_c_3_tile_v_5_3 = rf_matrix_c_3_tile_v_3_MPORT_5_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_3_tile_v_5_2 = rf_matrix_c_3_tile_v_2_MPORT_5_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_3_tile_v_5_1 = rf_matrix_c_3_tile_v_1_MPORT_5_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_3_tile_v_5_0 = rf_matrix_c_3_tile_v_0_MPORT_5_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_c_3_T_5 = {matrix_c_3_tile_v_5_3,matrix_c_3_tile_v_5_2,matrix_c_3_tile_v_5_1,
    matrix_c_3_tile_v_5_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [255:0] _GEN_4687 = 2'h3 == step ? _matrix_a_3_T_3 : matrix_a_3; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 159:21 212:23 247:27]
  wire [255:0] _GEN_4692 = 2'h3 == step ? _matrix_b_3_T_5 : matrix_b_3; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 160:21 212:23 248:27]
  wire [255:0] _GEN_4697 = 2'h3 == step ? _matrix_c_3_T_5 : matrix_c_3; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 161:21 212:23 249:27]
  wire [255:0] _GEN_4702 = 2'h2 == step ? _matrix_a_3_T_2 : _GEN_4687; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 212:23 241:27]
  wire [255:0] _GEN_4707 = 2'h2 == step ? _matrix_b_3_T_4 : _GEN_4692; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 212:23 242:27]
  wire [255:0] _GEN_4712 = 2'h2 == step ? _matrix_c_3_T_4 : _GEN_4697; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 212:23 243:27]
  wire [63:0] a_tile_v_78_1 = rf_a_tile_v_1_MPORT_78_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] a_tile_v_78_0 = rf_a_tile_v_0_MPORT_78_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_a_3_T_4 = {a_tile_v_78_1,a_tile_v_78_0,128'h0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 258:35]
  wire [63:0] matrix_b_3_tile_v_6_3 = rf_matrix_b_3_tile_v_3_MPORT_6_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_3_tile_v_6_2 = rf_matrix_b_3_tile_v_2_MPORT_6_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_3_tile_v_6_1 = rf_matrix_b_3_tile_v_1_MPORT_6_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_3_tile_v_6_0 = rf_matrix_b_3_tile_v_0_MPORT_6_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_b_3_T_6 = {matrix_b_3_tile_v_6_3,matrix_b_3_tile_v_6_2,matrix_b_3_tile_v_6_1,
    matrix_b_3_tile_v_6_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] matrix_c_3_tile_v_6_3 = rf_matrix_c_3_tile_v_3_MPORT_6_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_3_tile_v_6_2 = rf_matrix_c_3_tile_v_2_MPORT_6_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_3_tile_v_6_1 = rf_matrix_c_3_tile_v_1_MPORT_6_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_3_tile_v_6_0 = rf_matrix_c_3_tile_v_0_MPORT_6_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_c_3_T_6 = {matrix_c_3_tile_v_6_3,matrix_c_3_tile_v_6_2,matrix_c_3_tile_v_6_1,
    matrix_c_3_tile_v_6_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] a_tile_v_79_3 = rf_a_tile_v_3_MPORT_26_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] a_tile_v_79_2 = rf_a_tile_v_2_MPORT_26_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] a_tile_v_79_1 = rf_a_tile_v_1_MPORT_79_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] a_tile_v_79_0 = rf_a_tile_v_0_MPORT_79_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] a_79 = {a_tile_v_79_3,a_tile_v_79_2,a_tile_v_79_1,a_tile_v_79_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] matrix_b_3_tile_v_7_3 = rf_matrix_b_3_tile_v_3_MPORT_7_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_3_tile_v_7_2 = rf_matrix_b_3_tile_v_2_MPORT_7_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_3_tile_v_7_1 = rf_matrix_b_3_tile_v_1_MPORT_7_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_3_tile_v_7_0 = rf_matrix_b_3_tile_v_0_MPORT_7_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_b_3_T_7 = {matrix_b_3_tile_v_7_3,matrix_b_3_tile_v_7_2,matrix_b_3_tile_v_7_1,
    matrix_b_3_tile_v_7_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] matrix_c_3_tile_v_7_3 = rf_matrix_c_3_tile_v_3_MPORT_7_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_3_tile_v_7_2 = rf_matrix_c_3_tile_v_2_MPORT_7_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_3_tile_v_7_1 = rf_matrix_c_3_tile_v_1_MPORT_7_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_3_tile_v_7_0 = rf_matrix_c_3_tile_v_0_MPORT_7_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_c_3_T_7 = {matrix_c_3_tile_v_7_3,matrix_c_3_tile_v_7_2,matrix_c_3_tile_v_7_1,
    matrix_c_3_tile_v_7_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [255:0] _GEN_4857 = io_mixPc ? _matrix_a_3_T_4 : a_79; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 256:30 258:29 263:29]
  wire [255:0] _GEN_4858 = io_mixPc ? _matrix_b_3_T_6 : _matrix_b_3_T_7; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 256:30 259:29 264:29]
  wire [255:0] _GEN_4859 = io_mixPc ? _matrix_c_3_T_6 : _matrix_c_3_T_7; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 256:30 260:29 265:29]
  wire [63:0] a_tile_v_80_1 = rf_a_tile_v_1_MPORT_80_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] a_tile_v_80_0 = rf_a_tile_v_0_MPORT_80_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_a_3_T_5 = {a_tile_v_80_1,a_tile_v_80_0,128'h0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 271:35]
  wire [63:0] matrix_b_3_tile_v_8_3 = rf_matrix_b_3_tile_v_3_MPORT_8_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_3_tile_v_8_2 = rf_matrix_b_3_tile_v_2_MPORT_8_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_3_tile_v_8_1 = rf_matrix_b_3_tile_v_1_MPORT_8_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_3_tile_v_8_0 = rf_matrix_b_3_tile_v_0_MPORT_8_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_b_3_T_8 = {matrix_b_3_tile_v_8_3,matrix_b_3_tile_v_8_2,matrix_b_3_tile_v_8_1,
    matrix_b_3_tile_v_8_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] matrix_c_3_tile_v_8_3 = rf_matrix_c_3_tile_v_3_MPORT_8_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_3_tile_v_8_2 = rf_matrix_c_3_tile_v_2_MPORT_8_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_3_tile_v_8_1 = rf_matrix_c_3_tile_v_1_MPORT_8_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_3_tile_v_8_0 = rf_matrix_c_3_tile_v_0_MPORT_8_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_c_3_T_8 = {matrix_c_3_tile_v_8_3,matrix_c_3_tile_v_8_2,matrix_c_3_tile_v_8_1,
    matrix_c_3_tile_v_8_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] a_tile_v_81_3 = rf_a_tile_v_3_MPORT_27_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] a_tile_v_81_2 = rf_a_tile_v_2_MPORT_27_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] a_tile_v_81_1 = rf_a_tile_v_1_MPORT_81_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] a_tile_v_81_0 = rf_a_tile_v_0_MPORT_81_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] a_81 = {a_tile_v_81_3,a_tile_v_81_2,a_tile_v_81_1,a_tile_v_81_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] matrix_b_3_tile_v_9_3 = rf_matrix_b_3_tile_v_3_MPORT_9_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_3_tile_v_9_2 = rf_matrix_b_3_tile_v_2_MPORT_9_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_3_tile_v_9_1 = rf_matrix_b_3_tile_v_1_MPORT_9_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_3_tile_v_9_0 = rf_matrix_b_3_tile_v_0_MPORT_9_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_b_3_T_9 = {matrix_b_3_tile_v_9_3,matrix_b_3_tile_v_9_2,matrix_b_3_tile_v_9_1,
    matrix_b_3_tile_v_9_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] matrix_c_3_tile_v_9_3 = rf_matrix_c_3_tile_v_3_MPORT_9_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_3_tile_v_9_2 = rf_matrix_c_3_tile_v_2_MPORT_9_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_3_tile_v_9_1 = rf_matrix_c_3_tile_v_1_MPORT_9_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_3_tile_v_9_0 = rf_matrix_c_3_tile_v_0_MPORT_9_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_c_3_T_9 = {matrix_c_3_tile_v_9_3,matrix_c_3_tile_v_9_2,matrix_c_3_tile_v_9_1,
    matrix_c_3_tile_v_9_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [255:0] _GEN_4860 = io_mixPc ? _matrix_a_3_T_5 : a_81; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 269:30 271:29 276:29]
  wire [255:0] _GEN_4861 = io_mixPc ? _matrix_b_3_T_8 : _matrix_b_3_T_9; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 269:30 272:29 277:29]
  wire [255:0] _GEN_4862 = io_mixPc ? _matrix_c_3_T_8 : _matrix_c_3_T_9; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 269:30 273:29 278:29]
  wire [63:0] a_tile_v_82_1 = rf_a_tile_v_1_MPORT_82_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] a_tile_v_82_0 = rf_a_tile_v_0_MPORT_82_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_a_3_T_6 = {a_tile_v_82_1,a_tile_v_82_0,128'h0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 283:33]
  wire [63:0] matrix_b_3_tile_v_10_3 = rf_matrix_b_3_tile_v_3_MPORT_10_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_3_tile_v_10_2 = rf_matrix_b_3_tile_v_2_MPORT_10_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_3_tile_v_10_1 = rf_matrix_b_3_tile_v_1_MPORT_10_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_3_tile_v_10_0 = rf_matrix_b_3_tile_v_0_MPORT_10_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_b_3_T_10 = {matrix_b_3_tile_v_10_3,matrix_b_3_tile_v_10_2,matrix_b_3_tile_v_10_1,
    matrix_b_3_tile_v_10_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] matrix_c_3_tile_v_10_3 = rf_matrix_c_3_tile_v_3_MPORT_10_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_3_tile_v_10_2 = rf_matrix_c_3_tile_v_2_MPORT_10_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_3_tile_v_10_1 = rf_matrix_c_3_tile_v_1_MPORT_10_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_3_tile_v_10_0 = rf_matrix_c_3_tile_v_0_MPORT_10_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_c_3_T_10 = {matrix_c_3_tile_v_10_3,matrix_c_3_tile_v_10_2,matrix_c_3_tile_v_10_1,
    matrix_c_3_tile_v_10_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] a_tile_v_83_1 = rf_a_tile_v_1_MPORT_83_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] a_tile_v_83_0 = rf_a_tile_v_0_MPORT_83_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_a_3_T_7 = {a_tile_v_83_1,a_tile_v_83_0,128'h0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 289:33]
  wire [63:0] matrix_b_3_tile_v_11_3 = rf_matrix_b_3_tile_v_3_MPORT_11_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_3_tile_v_11_2 = rf_matrix_b_3_tile_v_2_MPORT_11_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_3_tile_v_11_1 = rf_matrix_b_3_tile_v_1_MPORT_11_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_3_tile_v_11_0 = rf_matrix_b_3_tile_v_0_MPORT_11_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_b_3_T_11 = {matrix_b_3_tile_v_11_3,matrix_b_3_tile_v_11_2,matrix_b_3_tile_v_11_1,
    matrix_b_3_tile_v_11_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] matrix_c_3_tile_v_11_3 = rf_matrix_c_3_tile_v_3_MPORT_11_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_3_tile_v_11_2 = rf_matrix_c_3_tile_v_2_MPORT_11_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_3_tile_v_11_1 = rf_matrix_c_3_tile_v_1_MPORT_11_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_3_tile_v_11_0 = rf_matrix_c_3_tile_v_0_MPORT_11_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_c_3_T_11 = {matrix_c_3_tile_v_11_3,matrix_c_3_tile_v_11_2,matrix_c_3_tile_v_11_1,
    matrix_c_3_tile_v_11_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [255:0] _GEN_4867 = _T_4 ? _matrix_a_3_T_7 : matrix_a_3; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 159:21 254:24 289:27]
  wire [255:0] _GEN_4872 = _T_4 ? _matrix_b_3_T_11 : matrix_b_3; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 160:21 254:24 290:27]
  wire [255:0] _GEN_4877 = _T_4 ? _matrix_c_3_T_11 : matrix_c_3; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 161:21 254:24 291:27]
  wire [255:0] _GEN_4882 = _T_3 ? _matrix_a_3_T_6 : _GEN_4867; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 254:24 283:27]
  wire [255:0] _GEN_4887 = _T_3 ? _matrix_b_3_T_10 : _GEN_4872; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 254:24 284:27]
  wire [255:0] _GEN_4892 = _T_3 ? _matrix_c_3_T_10 : _GEN_4877; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 254:24 285:27]
  wire [255:0] _GEN_4909 = _T_2 ? _GEN_4860 : _GEN_4882; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 254:24]
  wire [255:0] _GEN_4914 = _T_2 ? _GEN_4861 : _GEN_4887; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 254:24]
  wire [255:0] _GEN_4919 = _T_2 ? _GEN_4862 : _GEN_4892; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 254:24]
  wire [63:0] a_tile_v_84_1 = rf_a_tile_v_1_MPORT_84_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] a_tile_v_84_0 = rf_a_tile_v_0_MPORT_84_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_a_3_T_8 = {a_tile_v_84_1,a_tile_v_84_0,128'h0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 300:35]
  wire [63:0] matrix_b_3_tile_v_12_3 = rf_matrix_b_3_tile_v_3_MPORT_12_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_3_tile_v_12_2 = rf_matrix_b_3_tile_v_2_MPORT_12_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_3_tile_v_12_1 = rf_matrix_b_3_tile_v_1_MPORT_12_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_3_tile_v_12_0 = rf_matrix_b_3_tile_v_0_MPORT_12_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_b_3_T_12 = {matrix_b_3_tile_v_12_3,matrix_b_3_tile_v_12_2,matrix_b_3_tile_v_12_1,
    matrix_b_3_tile_v_12_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] matrix_c_3_tile_v_12_3 = rf_matrix_c_3_tile_v_3_MPORT_12_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_3_tile_v_12_2 = rf_matrix_c_3_tile_v_2_MPORT_12_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_3_tile_v_12_1 = rf_matrix_c_3_tile_v_1_MPORT_12_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_3_tile_v_12_0 = rf_matrix_c_3_tile_v_0_MPORT_12_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_c_3_T_12 = {matrix_c_3_tile_v_12_3,matrix_c_3_tile_v_12_2,matrix_c_3_tile_v_12_1,
    matrix_c_3_tile_v_12_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] a_tile_v_85_3 = rf_a_tile_v_3_MPORT_28_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] a_tile_v_85_2 = rf_a_tile_v_2_MPORT_28_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] a_tile_v_85_1 = rf_a_tile_v_1_MPORT_85_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] a_tile_v_85_0 = rf_a_tile_v_0_MPORT_85_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] a_85 = {a_tile_v_85_3,a_tile_v_85_2,a_tile_v_85_1,a_tile_v_85_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] matrix_b_3_tile_v_13_3 = rf_matrix_b_3_tile_v_3_MPORT_13_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_3_tile_v_13_2 = rf_matrix_b_3_tile_v_2_MPORT_13_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_3_tile_v_13_1 = rf_matrix_b_3_tile_v_1_MPORT_13_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_3_tile_v_13_0 = rf_matrix_b_3_tile_v_0_MPORT_13_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_b_3_T_13 = {matrix_b_3_tile_v_13_3,matrix_b_3_tile_v_13_2,matrix_b_3_tile_v_13_1,
    matrix_b_3_tile_v_13_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] matrix_c_3_tile_v_13_3 = rf_matrix_c_3_tile_v_3_MPORT_13_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_3_tile_v_13_2 = rf_matrix_c_3_tile_v_2_MPORT_13_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_3_tile_v_13_1 = rf_matrix_c_3_tile_v_1_MPORT_13_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_3_tile_v_13_0 = rf_matrix_c_3_tile_v_0_MPORT_13_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_c_3_T_13 = {matrix_c_3_tile_v_13_3,matrix_c_3_tile_v_13_2,matrix_c_3_tile_v_13_1,
    matrix_c_3_tile_v_13_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [255:0] _GEN_5037 = io_mixPc ? _matrix_a_3_T_8 : a_85; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 298:30 300:29 305:29]
  wire [255:0] _GEN_5038 = io_mixPc ? _matrix_b_3_T_12 : _matrix_b_3_T_13; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 298:30 301:29 306:29]
  wire [255:0] _GEN_5039 = io_mixPc ? _matrix_c_3_T_12 : _matrix_c_3_T_13; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 298:30 302:29 307:29]
  wire [63:0] a_tile_v_86_1 = rf_a_tile_v_1_MPORT_86_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] a_tile_v_86_0 = rf_a_tile_v_0_MPORT_86_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_a_3_T_9 = {a_tile_v_86_1,a_tile_v_86_0,128'h0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 313:35]
  wire [63:0] matrix_b_3_tile_v_14_3 = rf_matrix_b_3_tile_v_3_MPORT_14_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_3_tile_v_14_2 = rf_matrix_b_3_tile_v_2_MPORT_14_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_3_tile_v_14_1 = rf_matrix_b_3_tile_v_1_MPORT_14_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_3_tile_v_14_0 = rf_matrix_b_3_tile_v_0_MPORT_14_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_b_3_T_14 = {matrix_b_3_tile_v_14_3,matrix_b_3_tile_v_14_2,matrix_b_3_tile_v_14_1,
    matrix_b_3_tile_v_14_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] matrix_c_3_tile_v_14_3 = rf_matrix_c_3_tile_v_3_MPORT_14_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_3_tile_v_14_2 = rf_matrix_c_3_tile_v_2_MPORT_14_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_3_tile_v_14_1 = rf_matrix_c_3_tile_v_1_MPORT_14_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_3_tile_v_14_0 = rf_matrix_c_3_tile_v_0_MPORT_14_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_c_3_T_14 = {matrix_c_3_tile_v_14_3,matrix_c_3_tile_v_14_2,matrix_c_3_tile_v_14_1,
    matrix_c_3_tile_v_14_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] a_tile_v_87_3 = rf_a_tile_v_3_MPORT_29_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] a_tile_v_87_2 = rf_a_tile_v_2_MPORT_29_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] a_tile_v_87_1 = rf_a_tile_v_1_MPORT_87_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] a_tile_v_87_0 = rf_a_tile_v_0_MPORT_87_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] a_87 = {a_tile_v_87_3,a_tile_v_87_2,a_tile_v_87_1,a_tile_v_87_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] matrix_b_3_tile_v_15_3 = rf_matrix_b_3_tile_v_3_MPORT_15_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_3_tile_v_15_2 = rf_matrix_b_3_tile_v_2_MPORT_15_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_3_tile_v_15_1 = rf_matrix_b_3_tile_v_1_MPORT_15_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_3_tile_v_15_0 = rf_matrix_b_3_tile_v_0_MPORT_15_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_b_3_T_15 = {matrix_b_3_tile_v_15_3,matrix_b_3_tile_v_15_2,matrix_b_3_tile_v_15_1,
    matrix_b_3_tile_v_15_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] matrix_c_3_tile_v_15_3 = rf_matrix_c_3_tile_v_3_MPORT_15_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_3_tile_v_15_2 = rf_matrix_c_3_tile_v_2_MPORT_15_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_3_tile_v_15_1 = rf_matrix_c_3_tile_v_1_MPORT_15_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_3_tile_v_15_0 = rf_matrix_c_3_tile_v_0_MPORT_15_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_c_3_T_15 = {matrix_c_3_tile_v_15_3,matrix_c_3_tile_v_15_2,matrix_c_3_tile_v_15_1,
    matrix_c_3_tile_v_15_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [255:0] _GEN_5040 = io_mixPc ? _matrix_a_3_T_9 : a_87; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 311:30 313:29 318:29]
  wire [255:0] _GEN_5041 = io_mixPc ? _matrix_b_3_T_14 : _matrix_b_3_T_15; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 311:30 314:29 319:29]
  wire [255:0] _GEN_5042 = io_mixPc ? _matrix_c_3_T_14 : _matrix_c_3_T_15; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 311:30 315:29 320:29]
  wire [63:0] a_tile_v_88_1 = rf_a_tile_v_1_MPORT_88_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] a_tile_v_88_0 = rf_a_tile_v_0_MPORT_88_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_a_3_T_10 = {a_tile_v_88_1,a_tile_v_88_0,128'h0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 325:33]
  wire [63:0] matrix_b_3_tile_v_16_3 = rf_matrix_b_3_tile_v_3_MPORT_16_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_3_tile_v_16_2 = rf_matrix_b_3_tile_v_2_MPORT_16_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_3_tile_v_16_1 = rf_matrix_b_3_tile_v_1_MPORT_16_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_3_tile_v_16_0 = rf_matrix_b_3_tile_v_0_MPORT_16_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_b_3_T_16 = {matrix_b_3_tile_v_16_3,matrix_b_3_tile_v_16_2,matrix_b_3_tile_v_16_1,
    matrix_b_3_tile_v_16_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] matrix_c_3_tile_v_16_3 = rf_matrix_c_3_tile_v_3_MPORT_16_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_3_tile_v_16_2 = rf_matrix_c_3_tile_v_2_MPORT_16_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_3_tile_v_16_1 = rf_matrix_c_3_tile_v_1_MPORT_16_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_3_tile_v_16_0 = rf_matrix_c_3_tile_v_0_MPORT_16_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_c_3_T_16 = {matrix_c_3_tile_v_16_3,matrix_c_3_tile_v_16_2,matrix_c_3_tile_v_16_1,
    matrix_c_3_tile_v_16_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] a_tile_v_89_1 = rf_a_tile_v_1_MPORT_89_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] a_tile_v_89_0 = rf_a_tile_v_0_MPORT_89_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_a_3_T_11 = {a_tile_v_89_1,a_tile_v_89_0,128'h0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 331:33]
  wire [63:0] matrix_b_3_tile_v_17_3 = rf_matrix_b_3_tile_v_3_MPORT_17_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_3_tile_v_17_2 = rf_matrix_b_3_tile_v_2_MPORT_17_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_3_tile_v_17_1 = rf_matrix_b_3_tile_v_1_MPORT_17_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_3_tile_v_17_0 = rf_matrix_b_3_tile_v_0_MPORT_17_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_b_3_T_17 = {matrix_b_3_tile_v_17_3,matrix_b_3_tile_v_17_2,matrix_b_3_tile_v_17_1,
    matrix_b_3_tile_v_17_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] matrix_c_3_tile_v_17_3 = rf_matrix_c_3_tile_v_3_MPORT_17_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_3_tile_v_17_2 = rf_matrix_c_3_tile_v_2_MPORT_17_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_3_tile_v_17_1 = rf_matrix_c_3_tile_v_1_MPORT_17_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_3_tile_v_17_0 = rf_matrix_c_3_tile_v_0_MPORT_17_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_c_3_T_17 = {matrix_c_3_tile_v_17_3,matrix_c_3_tile_v_17_2,matrix_c_3_tile_v_17_1,
    matrix_c_3_tile_v_17_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [255:0] _GEN_5047 = _T_4 ? _matrix_a_3_T_11 : matrix_a_3; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 159:21 296:24 331:27]
  wire [255:0] _GEN_5052 = _T_4 ? _matrix_b_3_T_17 : matrix_b_3; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 160:21 296:24 332:27]
  wire [255:0] _GEN_5057 = _T_4 ? _matrix_c_3_T_17 : matrix_c_3; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 161:21 296:24 333:27]
  wire [255:0] _GEN_5062 = _T_3 ? _matrix_a_3_T_10 : _GEN_5047; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 296:24 325:27]
  wire [255:0] _GEN_5067 = _T_3 ? _matrix_b_3_T_16 : _GEN_5052; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 296:24 326:27]
  wire [255:0] _GEN_5072 = _T_3 ? _matrix_c_3_T_16 : _GEN_5057; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 296:24 327:27]
  wire [255:0] _GEN_5089 = _T_2 ? _GEN_5040 : _GEN_5062; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 296:24]
  wire [255:0] _GEN_5094 = _T_2 ? _GEN_5041 : _GEN_5067; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 296:24]
  wire [255:0] _GEN_5099 = _T_2 ? _GEN_5042 : _GEN_5072; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 296:24]
  wire [255:0] _GEN_5142 = _T_1 ? _GEN_5037 : _GEN_5089; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 296:24]
  wire [255:0] _GEN_5147 = _T_1 ? _GEN_5038 : _GEN_5094; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 296:24]
  wire [255:0] _GEN_5152 = _T_1 ? _GEN_5039 : _GEN_5099; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 296:24]
  wire [63:0] a_tile_v_90_1 = rf_a_tile_v_1_MPORT_90_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] a_tile_v_90_0 = rf_a_tile_v_0_MPORT_90_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_a_3_T_12 = {a_tile_v_90_1,a_tile_v_90_0,128'h0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 342:35]
  wire [63:0] matrix_b_3_tile_v_18_3 = rf_matrix_b_3_tile_v_3_MPORT_18_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_3_tile_v_18_2 = rf_matrix_b_3_tile_v_2_MPORT_18_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_3_tile_v_18_1 = rf_matrix_b_3_tile_v_1_MPORT_18_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_3_tile_v_18_0 = rf_matrix_b_3_tile_v_0_MPORT_18_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_b_3_T_18 = {matrix_b_3_tile_v_18_3,matrix_b_3_tile_v_18_2,matrix_b_3_tile_v_18_1,
    matrix_b_3_tile_v_18_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] matrix_c_3_tile_v_18_3 = rf_matrix_c_3_tile_v_3_MPORT_18_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_3_tile_v_18_2 = rf_matrix_c_3_tile_v_2_MPORT_18_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_3_tile_v_18_1 = rf_matrix_c_3_tile_v_1_MPORT_18_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_3_tile_v_18_0 = rf_matrix_c_3_tile_v_0_MPORT_18_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_c_3_T_18 = {matrix_c_3_tile_v_18_3,matrix_c_3_tile_v_18_2,matrix_c_3_tile_v_18_1,
    matrix_c_3_tile_v_18_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] a_tile_v_91_3 = rf_a_tile_v_3_MPORT_30_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] a_tile_v_91_2 = rf_a_tile_v_2_MPORT_30_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] a_tile_v_91_1 = rf_a_tile_v_1_MPORT_91_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] a_tile_v_91_0 = rf_a_tile_v_0_MPORT_91_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] a_91 = {a_tile_v_91_3,a_tile_v_91_2,a_tile_v_91_1,a_tile_v_91_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] matrix_b_3_tile_v_19_3 = rf_matrix_b_3_tile_v_3_MPORT_19_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_3_tile_v_19_2 = rf_matrix_b_3_tile_v_2_MPORT_19_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_3_tile_v_19_1 = rf_matrix_b_3_tile_v_1_MPORT_19_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_3_tile_v_19_0 = rf_matrix_b_3_tile_v_0_MPORT_19_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_b_3_T_19 = {matrix_b_3_tile_v_19_3,matrix_b_3_tile_v_19_2,matrix_b_3_tile_v_19_1,
    matrix_b_3_tile_v_19_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] matrix_c_3_tile_v_19_3 = rf_matrix_c_3_tile_v_3_MPORT_19_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_3_tile_v_19_2 = rf_matrix_c_3_tile_v_2_MPORT_19_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_3_tile_v_19_1 = rf_matrix_c_3_tile_v_1_MPORT_19_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_3_tile_v_19_0 = rf_matrix_c_3_tile_v_0_MPORT_19_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_c_3_T_19 = {matrix_c_3_tile_v_19_3,matrix_c_3_tile_v_19_2,matrix_c_3_tile_v_19_1,
    matrix_c_3_tile_v_19_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [255:0] _GEN_5217 = io_mixPc ? _matrix_a_3_T_12 : a_91; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 340:30 342:29 347:29]
  wire [255:0] _GEN_5218 = io_mixPc ? _matrix_b_3_T_18 : _matrix_b_3_T_19; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 340:30 343:29 348:29]
  wire [255:0] _GEN_5219 = io_mixPc ? _matrix_c_3_T_18 : _matrix_c_3_T_19; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 340:30 344:29 349:29]
  wire [63:0] a_tile_v_92_1 = rf_a_tile_v_1_MPORT_92_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] a_tile_v_92_0 = rf_a_tile_v_0_MPORT_92_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_a_3_T_13 = {a_tile_v_92_1,a_tile_v_92_0,128'h0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 355:35]
  wire [63:0] matrix_b_3_tile_v_20_3 = rf_matrix_b_3_tile_v_3_MPORT_20_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_3_tile_v_20_2 = rf_matrix_b_3_tile_v_2_MPORT_20_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_3_tile_v_20_1 = rf_matrix_b_3_tile_v_1_MPORT_20_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_3_tile_v_20_0 = rf_matrix_b_3_tile_v_0_MPORT_20_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_b_3_T_20 = {matrix_b_3_tile_v_20_3,matrix_b_3_tile_v_20_2,matrix_b_3_tile_v_20_1,
    matrix_b_3_tile_v_20_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] matrix_c_3_tile_v_20_3 = rf_matrix_c_3_tile_v_3_MPORT_20_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_3_tile_v_20_2 = rf_matrix_c_3_tile_v_2_MPORT_20_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_3_tile_v_20_1 = rf_matrix_c_3_tile_v_1_MPORT_20_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_3_tile_v_20_0 = rf_matrix_c_3_tile_v_0_MPORT_20_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_c_3_T_20 = {matrix_c_3_tile_v_20_3,matrix_c_3_tile_v_20_2,matrix_c_3_tile_v_20_1,
    matrix_c_3_tile_v_20_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] a_tile_v_93_3 = rf_a_tile_v_3_MPORT_31_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] a_tile_v_93_2 = rf_a_tile_v_2_MPORT_31_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] a_tile_v_93_1 = rf_a_tile_v_1_MPORT_93_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] a_tile_v_93_0 = rf_a_tile_v_0_MPORT_93_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] a_93 = {a_tile_v_93_3,a_tile_v_93_2,a_tile_v_93_1,a_tile_v_93_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] matrix_b_3_tile_v_21_3 = rf_matrix_b_3_tile_v_3_MPORT_21_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_3_tile_v_21_2 = rf_matrix_b_3_tile_v_2_MPORT_21_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_3_tile_v_21_1 = rf_matrix_b_3_tile_v_1_MPORT_21_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_3_tile_v_21_0 = rf_matrix_b_3_tile_v_0_MPORT_21_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_b_3_T_21 = {matrix_b_3_tile_v_21_3,matrix_b_3_tile_v_21_2,matrix_b_3_tile_v_21_1,
    matrix_b_3_tile_v_21_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] matrix_c_3_tile_v_21_3 = rf_matrix_c_3_tile_v_3_MPORT_21_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_3_tile_v_21_2 = rf_matrix_c_3_tile_v_2_MPORT_21_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_3_tile_v_21_1 = rf_matrix_c_3_tile_v_1_MPORT_21_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_3_tile_v_21_0 = rf_matrix_c_3_tile_v_0_MPORT_21_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_c_3_T_21 = {matrix_c_3_tile_v_21_3,matrix_c_3_tile_v_21_2,matrix_c_3_tile_v_21_1,
    matrix_c_3_tile_v_21_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [255:0] _GEN_5220 = io_mixPc ? _matrix_a_3_T_13 : a_93; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 353:30 355:29 360:29]
  wire [255:0] _GEN_5221 = io_mixPc ? _matrix_b_3_T_20 : _matrix_b_3_T_21; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 353:30 356:29 361:29]
  wire [255:0] _GEN_5222 = io_mixPc ? _matrix_c_3_T_20 : _matrix_c_3_T_21; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 353:30 357:29 362:29]
  wire [63:0] a_tile_v_94_1 = rf_a_tile_v_1_MPORT_94_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] a_tile_v_94_0 = rf_a_tile_v_0_MPORT_94_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_a_3_T_14 = {a_tile_v_94_1,a_tile_v_94_0,128'h0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 367:33]
  wire [63:0] matrix_b_3_tile_v_22_3 = rf_matrix_b_3_tile_v_3_MPORT_22_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_3_tile_v_22_2 = rf_matrix_b_3_tile_v_2_MPORT_22_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_3_tile_v_22_1 = rf_matrix_b_3_tile_v_1_MPORT_22_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_3_tile_v_22_0 = rf_matrix_b_3_tile_v_0_MPORT_22_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_b_3_T_22 = {matrix_b_3_tile_v_22_3,matrix_b_3_tile_v_22_2,matrix_b_3_tile_v_22_1,
    matrix_b_3_tile_v_22_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] matrix_c_3_tile_v_22_3 = rf_matrix_c_3_tile_v_3_MPORT_22_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_3_tile_v_22_2 = rf_matrix_c_3_tile_v_2_MPORT_22_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_3_tile_v_22_1 = rf_matrix_c_3_tile_v_1_MPORT_22_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_3_tile_v_22_0 = rf_matrix_c_3_tile_v_0_MPORT_22_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_c_3_T_22 = {matrix_c_3_tile_v_22_3,matrix_c_3_tile_v_22_2,matrix_c_3_tile_v_22_1,
    matrix_c_3_tile_v_22_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] a_tile_v_95_1 = rf_a_tile_v_1_MPORT_95_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] a_tile_v_95_0 = rf_a_tile_v_0_MPORT_95_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_a_3_T_15 = {a_tile_v_95_1,a_tile_v_95_0,128'h0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 373:33]
  wire [63:0] matrix_b_3_tile_v_23_3 = rf_matrix_b_3_tile_v_3_MPORT_23_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_3_tile_v_23_2 = rf_matrix_b_3_tile_v_2_MPORT_23_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_3_tile_v_23_1 = rf_matrix_b_3_tile_v_1_MPORT_23_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_3_tile_v_23_0 = rf_matrix_b_3_tile_v_0_MPORT_23_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_b_3_T_23 = {matrix_b_3_tile_v_23_3,matrix_b_3_tile_v_23_2,matrix_b_3_tile_v_23_1,
    matrix_b_3_tile_v_23_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] matrix_c_3_tile_v_23_3 = rf_matrix_c_3_tile_v_3_MPORT_23_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_3_tile_v_23_2 = rf_matrix_c_3_tile_v_2_MPORT_23_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_3_tile_v_23_1 = rf_matrix_c_3_tile_v_1_MPORT_23_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_3_tile_v_23_0 = rf_matrix_c_3_tile_v_0_MPORT_23_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_c_3_T_23 = {matrix_c_3_tile_v_23_3,matrix_c_3_tile_v_23_2,matrix_c_3_tile_v_23_1,
    matrix_c_3_tile_v_23_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [255:0] _GEN_5227 = _T_4 ? _matrix_a_3_T_15 : matrix_a_3; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 159:21 338:24 373:27]
  wire [255:0] _GEN_5232 = _T_4 ? _matrix_b_3_T_23 : matrix_b_3; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 160:21 338:24 374:27]
  wire [255:0] _GEN_5237 = _T_4 ? _matrix_c_3_T_23 : matrix_c_3; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 161:21 338:24 375:27]
  wire [255:0] _GEN_5242 = _T_3 ? _matrix_a_3_T_14 : _GEN_5227; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 338:24 367:27]
  wire [255:0] _GEN_5247 = _T_3 ? _matrix_b_3_T_22 : _GEN_5232; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 338:24 368:27]
  wire [255:0] _GEN_5252 = _T_3 ? _matrix_c_3_T_22 : _GEN_5237; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 338:24 369:27]
  wire [255:0] _GEN_5269 = _T_2 ? _GEN_5220 : _GEN_5242; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 338:24]
  wire [255:0] _GEN_5274 = _T_2 ? _GEN_5221 : _GEN_5247; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 338:24]
  wire [255:0] _GEN_5279 = _T_2 ? _GEN_5222 : _GEN_5252; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 338:24]
  wire [255:0] _GEN_5322 = _T_1 ? _GEN_5217 : _GEN_5269; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 338:24]
  wire [255:0] _GEN_5327 = _T_1 ? _GEN_5218 : _GEN_5274; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 338:24]
  wire [255:0] _GEN_5332 = _T_1 ? _GEN_5219 : _GEN_5279; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 338:24]
  wire [255:0] _GEN_5401 = 2'h3 == set ? _GEN_5322 : matrix_a_3; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 210:18 159:21]
  wire [255:0] _GEN_5406 = 2'h3 == set ? _GEN_5327 : matrix_b_3; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 210:18 160:21]
  wire [255:0] _GEN_5411 = 2'h3 == set ? _GEN_5332 : matrix_c_3; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 210:18 161:21]
  wire [63:0] a_tile_v_96_1 = rf_a_tile_v_1_MPORT_96_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] a_tile_v_96_0 = rf_a_tile_v_0_MPORT_96_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_a_4_T = {a_tile_v_96_1,a_tile_v_96_0,128'h0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 216:35]
  wire [63:0] matrix_b_4_tile_v__3 = rf_matrix_b_4_tile_v_3_MPORT_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_4_tile_v__2 = rf_matrix_b_4_tile_v_2_MPORT_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_4_tile_v__1 = rf_matrix_b_4_tile_v_1_MPORT_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_4_tile_v__0 = rf_matrix_b_4_tile_v_0_MPORT_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_b_4_T = {matrix_b_4_tile_v__3,matrix_b_4_tile_v__2,matrix_b_4_tile_v__1,matrix_b_4_tile_v__0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] matrix_c_4_tile_v__3 = rf_matrix_c_4_tile_v_3_MPORT_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_4_tile_v__2 = rf_matrix_c_4_tile_v_2_MPORT_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_4_tile_v__1 = rf_matrix_c_4_tile_v_1_MPORT_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_4_tile_v__0 = rf_matrix_c_4_tile_v_0_MPORT_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_c_4_T = {matrix_c_4_tile_v__3,matrix_c_4_tile_v__2,matrix_c_4_tile_v__1,matrix_c_4_tile_v__0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] a_tile_v_97_3 = rf_a_tile_v_3_MPORT_32_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] a_tile_v_97_2 = rf_a_tile_v_2_MPORT_32_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] a_tile_v_97_1 = rf_a_tile_v_1_MPORT_97_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] a_tile_v_97_0 = rf_a_tile_v_0_MPORT_97_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] a_97 = {a_tile_v_97_3,a_tile_v_97_2,a_tile_v_97_1,a_tile_v_97_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] matrix_b_4_tile_v_1_3 = rf_matrix_b_4_tile_v_3_MPORT_1_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_4_tile_v_1_2 = rf_matrix_b_4_tile_v_2_MPORT_1_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_4_tile_v_1_1 = rf_matrix_b_4_tile_v_1_MPORT_1_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_4_tile_v_1_0 = rf_matrix_b_4_tile_v_0_MPORT_1_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_b_4_T_1 = {matrix_b_4_tile_v_1_3,matrix_b_4_tile_v_1_2,matrix_b_4_tile_v_1_1,
    matrix_b_4_tile_v_1_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] matrix_c_4_tile_v_1_3 = rf_matrix_c_4_tile_v_3_MPORT_1_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_4_tile_v_1_2 = rf_matrix_c_4_tile_v_2_MPORT_1_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_4_tile_v_1_1 = rf_matrix_c_4_tile_v_1_MPORT_1_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_4_tile_v_1_0 = rf_matrix_c_4_tile_v_0_MPORT_1_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_c_4_T_1 = {matrix_c_4_tile_v_1_3,matrix_c_4_tile_v_1_2,matrix_c_4_tile_v_1_1,
    matrix_c_4_tile_v_1_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] a_tile_v_98_1 = rf_a_tile_v_1_MPORT_98_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] a_tile_v_98_0 = rf_a_tile_v_0_MPORT_98_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_a_4_T_1 = {a_tile_v_98_1,a_tile_v_98_0,128'h0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 229:35]
  wire [63:0] matrix_b_4_tile_v_2_3 = rf_matrix_b_4_tile_v_3_MPORT_2_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_4_tile_v_2_2 = rf_matrix_b_4_tile_v_2_MPORT_2_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_4_tile_v_2_1 = rf_matrix_b_4_tile_v_1_MPORT_2_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_4_tile_v_2_0 = rf_matrix_b_4_tile_v_0_MPORT_2_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_b_4_T_2 = {matrix_b_4_tile_v_2_3,matrix_b_4_tile_v_2_2,matrix_b_4_tile_v_2_1,
    matrix_b_4_tile_v_2_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] matrix_c_4_tile_v_2_3 = rf_matrix_c_4_tile_v_3_MPORT_2_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_4_tile_v_2_2 = rf_matrix_c_4_tile_v_2_MPORT_2_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_4_tile_v_2_1 = rf_matrix_c_4_tile_v_1_MPORT_2_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_4_tile_v_2_0 = rf_matrix_c_4_tile_v_0_MPORT_2_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_c_4_T_2 = {matrix_c_4_tile_v_2_3,matrix_c_4_tile_v_2_2,matrix_c_4_tile_v_2_1,
    matrix_c_4_tile_v_2_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] a_tile_v_99_3 = rf_a_tile_v_3_MPORT_33_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] a_tile_v_99_2 = rf_a_tile_v_2_MPORT_33_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] a_tile_v_99_1 = rf_a_tile_v_1_MPORT_99_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] a_tile_v_99_0 = rf_a_tile_v_0_MPORT_99_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] a_99 = {a_tile_v_99_3,a_tile_v_99_2,a_tile_v_99_1,a_tile_v_99_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] matrix_b_4_tile_v_3_3 = rf_matrix_b_4_tile_v_3_MPORT_3_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_4_tile_v_3_2 = rf_matrix_b_4_tile_v_2_MPORT_3_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_4_tile_v_3_1 = rf_matrix_b_4_tile_v_1_MPORT_3_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_4_tile_v_3_0 = rf_matrix_b_4_tile_v_0_MPORT_3_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_b_4_T_3 = {matrix_b_4_tile_v_3_3,matrix_b_4_tile_v_3_2,matrix_b_4_tile_v_3_1,
    matrix_b_4_tile_v_3_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] matrix_c_4_tile_v_3_3 = rf_matrix_c_4_tile_v_3_MPORT_3_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_4_tile_v_3_2 = rf_matrix_c_4_tile_v_2_MPORT_3_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_4_tile_v_3_1 = rf_matrix_c_4_tile_v_1_MPORT_3_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_4_tile_v_3_0 = rf_matrix_c_4_tile_v_0_MPORT_3_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_c_4_T_3 = {matrix_c_4_tile_v_3_3,matrix_c_4_tile_v_3_2,matrix_c_4_tile_v_3_1,
    matrix_c_4_tile_v_3_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [255:0] _GEN_6196 = io_mixPc ? _matrix_a_4_T_1 : a_99; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 227:30 229:29 234:29]
  wire [255:0] _GEN_6197 = io_mixPc ? _matrix_b_4_T_2 : _matrix_b_4_T_3; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 227:30 230:29 235:29]
  wire [255:0] _GEN_6202 = io_mixPc ? _matrix_c_4_T_2 : _matrix_c_4_T_3; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 227:30 231:29 236:29]
  wire [63:0] a_tile_v_100_1 = rf_a_tile_v_1_MPORT_100_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] a_tile_v_100_0 = rf_a_tile_v_0_MPORT_100_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_a_4_T_2 = {a_tile_v_100_1,a_tile_v_100_0,128'h0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 241:33]
  wire [63:0] matrix_b_4_tile_v_4_3 = rf_matrix_b_4_tile_v_3_MPORT_4_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_4_tile_v_4_2 = rf_matrix_b_4_tile_v_2_MPORT_4_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_4_tile_v_4_1 = rf_matrix_b_4_tile_v_1_MPORT_4_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_4_tile_v_4_0 = rf_matrix_b_4_tile_v_0_MPORT_4_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_b_4_T_4 = {matrix_b_4_tile_v_4_3,matrix_b_4_tile_v_4_2,matrix_b_4_tile_v_4_1,
    matrix_b_4_tile_v_4_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] matrix_c_4_tile_v_4_3 = rf_matrix_c_4_tile_v_3_MPORT_4_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_4_tile_v_4_2 = rf_matrix_c_4_tile_v_2_MPORT_4_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_4_tile_v_4_1 = rf_matrix_c_4_tile_v_1_MPORT_4_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_4_tile_v_4_0 = rf_matrix_c_4_tile_v_0_MPORT_4_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_c_4_T_4 = {matrix_c_4_tile_v_4_3,matrix_c_4_tile_v_4_2,matrix_c_4_tile_v_4_1,
    matrix_c_4_tile_v_4_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] a_tile_v_101_1 = rf_a_tile_v_1_MPORT_101_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] a_tile_v_101_0 = rf_a_tile_v_0_MPORT_101_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_a_4_T_3 = {a_tile_v_101_1,a_tile_v_101_0,128'h0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 247:33]
  wire [63:0] matrix_b_4_tile_v_5_3 = rf_matrix_b_4_tile_v_3_MPORT_5_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_4_tile_v_5_2 = rf_matrix_b_4_tile_v_2_MPORT_5_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_4_tile_v_5_1 = rf_matrix_b_4_tile_v_1_MPORT_5_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_4_tile_v_5_0 = rf_matrix_b_4_tile_v_0_MPORT_5_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_b_4_T_5 = {matrix_b_4_tile_v_5_3,matrix_b_4_tile_v_5_2,matrix_b_4_tile_v_5_1,
    matrix_b_4_tile_v_5_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] matrix_c_4_tile_v_5_3 = rf_matrix_c_4_tile_v_3_MPORT_5_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_4_tile_v_5_2 = rf_matrix_c_4_tile_v_2_MPORT_5_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_4_tile_v_5_1 = rf_matrix_c_4_tile_v_1_MPORT_5_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_4_tile_v_5_0 = rf_matrix_c_4_tile_v_0_MPORT_5_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_c_4_T_5 = {matrix_c_4_tile_v_5_3,matrix_c_4_tile_v_5_2,matrix_c_4_tile_v_5_1,
    matrix_c_4_tile_v_5_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [255:0] _GEN_6211 = 2'h3 == step ? _matrix_a_4_T_3 : matrix_a_4; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 159:21 212:23 247:27]
  wire [255:0] _GEN_6216 = 2'h3 == step ? _matrix_b_4_T_5 : matrix_b_4; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 160:21 212:23 248:27]
  wire [255:0] _GEN_6221 = 2'h3 == step ? _matrix_c_4_T_5 : matrix_c_4; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 161:21 212:23 249:27]
  wire [255:0] _GEN_6226 = 2'h2 == step ? _matrix_a_4_T_2 : _GEN_6211; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 212:23 241:27]
  wire [255:0] _GEN_6231 = 2'h2 == step ? _matrix_b_4_T_4 : _GEN_6216; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 212:23 242:27]
  wire [255:0] _GEN_6236 = 2'h2 == step ? _matrix_c_4_T_4 : _GEN_6221; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 212:23 243:27]
  wire [63:0] a_tile_v_102_1 = rf_a_tile_v_1_MPORT_102_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] a_tile_v_102_0 = rf_a_tile_v_0_MPORT_102_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_a_4_T_4 = {a_tile_v_102_1,a_tile_v_102_0,128'h0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 258:35]
  wire [63:0] matrix_b_4_tile_v_6_3 = rf_matrix_b_4_tile_v_3_MPORT_6_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_4_tile_v_6_2 = rf_matrix_b_4_tile_v_2_MPORT_6_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_4_tile_v_6_1 = rf_matrix_b_4_tile_v_1_MPORT_6_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_4_tile_v_6_0 = rf_matrix_b_4_tile_v_0_MPORT_6_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_b_4_T_6 = {matrix_b_4_tile_v_6_3,matrix_b_4_tile_v_6_2,matrix_b_4_tile_v_6_1,
    matrix_b_4_tile_v_6_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] matrix_c_4_tile_v_6_3 = rf_matrix_c_4_tile_v_3_MPORT_6_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_4_tile_v_6_2 = rf_matrix_c_4_tile_v_2_MPORT_6_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_4_tile_v_6_1 = rf_matrix_c_4_tile_v_1_MPORT_6_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_4_tile_v_6_0 = rf_matrix_c_4_tile_v_0_MPORT_6_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_c_4_T_6 = {matrix_c_4_tile_v_6_3,matrix_c_4_tile_v_6_2,matrix_c_4_tile_v_6_1,
    matrix_c_4_tile_v_6_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] a_tile_v_103_3 = rf_a_tile_v_3_MPORT_34_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] a_tile_v_103_2 = rf_a_tile_v_2_MPORT_34_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] a_tile_v_103_1 = rf_a_tile_v_1_MPORT_103_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] a_tile_v_103_0 = rf_a_tile_v_0_MPORT_103_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] a_103 = {a_tile_v_103_3,a_tile_v_103_2,a_tile_v_103_1,a_tile_v_103_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] matrix_b_4_tile_v_7_3 = rf_matrix_b_4_tile_v_3_MPORT_7_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_4_tile_v_7_2 = rf_matrix_b_4_tile_v_2_MPORT_7_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_4_tile_v_7_1 = rf_matrix_b_4_tile_v_1_MPORT_7_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_4_tile_v_7_0 = rf_matrix_b_4_tile_v_0_MPORT_7_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_b_4_T_7 = {matrix_b_4_tile_v_7_3,matrix_b_4_tile_v_7_2,matrix_b_4_tile_v_7_1,
    matrix_b_4_tile_v_7_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] matrix_c_4_tile_v_7_3 = rf_matrix_c_4_tile_v_3_MPORT_7_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_4_tile_v_7_2 = rf_matrix_c_4_tile_v_2_MPORT_7_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_4_tile_v_7_1 = rf_matrix_c_4_tile_v_1_MPORT_7_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_4_tile_v_7_0 = rf_matrix_c_4_tile_v_0_MPORT_7_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_c_4_T_7 = {matrix_c_4_tile_v_7_3,matrix_c_4_tile_v_7_2,matrix_c_4_tile_v_7_1,
    matrix_c_4_tile_v_7_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [255:0] _GEN_6383 = io_mixPc ? _matrix_a_4_T_4 : a_103; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 256:30 258:29 263:29]
  wire [255:0] _GEN_6388 = io_mixPc ? _matrix_b_4_T_6 : _matrix_b_4_T_7; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 256:30 259:29 264:29]
  wire [255:0] _GEN_6389 = io_mixPc ? _matrix_c_4_T_6 : _matrix_c_4_T_7; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 256:30 260:29 265:29]
  wire [63:0] a_tile_v_104_1 = rf_a_tile_v_1_MPORT_104_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] a_tile_v_104_0 = rf_a_tile_v_0_MPORT_104_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_a_4_T_5 = {a_tile_v_104_1,a_tile_v_104_0,128'h0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 271:35]
  wire [63:0] matrix_b_4_tile_v_8_3 = rf_matrix_b_4_tile_v_3_MPORT_8_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_4_tile_v_8_2 = rf_matrix_b_4_tile_v_2_MPORT_8_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_4_tile_v_8_1 = rf_matrix_b_4_tile_v_1_MPORT_8_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_4_tile_v_8_0 = rf_matrix_b_4_tile_v_0_MPORT_8_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_b_4_T_8 = {matrix_b_4_tile_v_8_3,matrix_b_4_tile_v_8_2,matrix_b_4_tile_v_8_1,
    matrix_b_4_tile_v_8_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] matrix_c_4_tile_v_8_3 = rf_matrix_c_4_tile_v_3_MPORT_8_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_4_tile_v_8_2 = rf_matrix_c_4_tile_v_2_MPORT_8_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_4_tile_v_8_1 = rf_matrix_c_4_tile_v_1_MPORT_8_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_4_tile_v_8_0 = rf_matrix_c_4_tile_v_0_MPORT_8_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_c_4_T_8 = {matrix_c_4_tile_v_8_3,matrix_c_4_tile_v_8_2,matrix_c_4_tile_v_8_1,
    matrix_c_4_tile_v_8_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] a_tile_v_105_3 = rf_a_tile_v_3_MPORT_35_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] a_tile_v_105_2 = rf_a_tile_v_2_MPORT_35_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] a_tile_v_105_1 = rf_a_tile_v_1_MPORT_105_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] a_tile_v_105_0 = rf_a_tile_v_0_MPORT_105_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] a_105 = {a_tile_v_105_3,a_tile_v_105_2,a_tile_v_105_1,a_tile_v_105_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] matrix_b_4_tile_v_9_3 = rf_matrix_b_4_tile_v_3_MPORT_9_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_4_tile_v_9_2 = rf_matrix_b_4_tile_v_2_MPORT_9_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_4_tile_v_9_1 = rf_matrix_b_4_tile_v_1_MPORT_9_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_4_tile_v_9_0 = rf_matrix_b_4_tile_v_0_MPORT_9_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_b_4_T_9 = {matrix_b_4_tile_v_9_3,matrix_b_4_tile_v_9_2,matrix_b_4_tile_v_9_1,
    matrix_b_4_tile_v_9_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] matrix_c_4_tile_v_9_3 = rf_matrix_c_4_tile_v_3_MPORT_9_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_4_tile_v_9_2 = rf_matrix_c_4_tile_v_2_MPORT_9_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_4_tile_v_9_1 = rf_matrix_c_4_tile_v_1_MPORT_9_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_4_tile_v_9_0 = rf_matrix_c_4_tile_v_0_MPORT_9_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_c_4_T_9 = {matrix_c_4_tile_v_9_3,matrix_c_4_tile_v_9_2,matrix_c_4_tile_v_9_1,
    matrix_c_4_tile_v_9_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [255:0] _GEN_6400 = io_mixPc ? _matrix_a_4_T_5 : a_105; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 269:30 271:29 276:29]
  wire [255:0] _GEN_6401 = io_mixPc ? _matrix_b_4_T_8 : _matrix_b_4_T_9; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 269:30 272:29 277:29]
  wire [255:0] _GEN_6402 = io_mixPc ? _matrix_c_4_T_8 : _matrix_c_4_T_9; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 269:30 273:29 278:29]
  wire [63:0] a_tile_v_106_1 = rf_a_tile_v_1_MPORT_106_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] a_tile_v_106_0 = rf_a_tile_v_0_MPORT_106_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_a_4_T_6 = {a_tile_v_106_1,a_tile_v_106_0,128'h0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 283:33]
  wire [63:0] matrix_b_4_tile_v_10_3 = rf_matrix_b_4_tile_v_3_MPORT_10_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_4_tile_v_10_2 = rf_matrix_b_4_tile_v_2_MPORT_10_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_4_tile_v_10_1 = rf_matrix_b_4_tile_v_1_MPORT_10_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_4_tile_v_10_0 = rf_matrix_b_4_tile_v_0_MPORT_10_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_b_4_T_10 = {matrix_b_4_tile_v_10_3,matrix_b_4_tile_v_10_2,matrix_b_4_tile_v_10_1,
    matrix_b_4_tile_v_10_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] matrix_c_4_tile_v_10_3 = rf_matrix_c_4_tile_v_3_MPORT_10_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_4_tile_v_10_2 = rf_matrix_c_4_tile_v_2_MPORT_10_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_4_tile_v_10_1 = rf_matrix_c_4_tile_v_1_MPORT_10_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_4_tile_v_10_0 = rf_matrix_c_4_tile_v_0_MPORT_10_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_c_4_T_10 = {matrix_c_4_tile_v_10_3,matrix_c_4_tile_v_10_2,matrix_c_4_tile_v_10_1,
    matrix_c_4_tile_v_10_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] a_tile_v_107_1 = rf_a_tile_v_1_MPORT_107_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] a_tile_v_107_0 = rf_a_tile_v_0_MPORT_107_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_a_4_T_7 = {a_tile_v_107_1,a_tile_v_107_0,128'h0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 289:33]
  wire [63:0] matrix_b_4_tile_v_11_3 = rf_matrix_b_4_tile_v_3_MPORT_11_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_4_tile_v_11_2 = rf_matrix_b_4_tile_v_2_MPORT_11_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_4_tile_v_11_1 = rf_matrix_b_4_tile_v_1_MPORT_11_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_4_tile_v_11_0 = rf_matrix_b_4_tile_v_0_MPORT_11_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_b_4_T_11 = {matrix_b_4_tile_v_11_3,matrix_b_4_tile_v_11_2,matrix_b_4_tile_v_11_1,
    matrix_b_4_tile_v_11_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] matrix_c_4_tile_v_11_3 = rf_matrix_c_4_tile_v_3_MPORT_11_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_4_tile_v_11_2 = rf_matrix_c_4_tile_v_2_MPORT_11_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_4_tile_v_11_1 = rf_matrix_c_4_tile_v_1_MPORT_11_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_4_tile_v_11_0 = rf_matrix_c_4_tile_v_0_MPORT_11_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_c_4_T_11 = {matrix_c_4_tile_v_11_3,matrix_c_4_tile_v_11_2,matrix_c_4_tile_v_11_1,
    matrix_c_4_tile_v_11_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [255:0] _GEN_6407 = _T_4 ? _matrix_a_4_T_7 : matrix_a_4; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 159:21 254:24 289:27]
  wire [255:0] _GEN_6412 = _T_4 ? _matrix_b_4_T_11 : matrix_b_4; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 160:21 254:24 290:27]
  wire [255:0] _GEN_6417 = _T_4 ? _matrix_c_4_T_11 : matrix_c_4; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 161:21 254:24 291:27]
  wire [255:0] _GEN_6422 = _T_3 ? _matrix_a_4_T_6 : _GEN_6407; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 254:24 283:27]
  wire [255:0] _GEN_6427 = _T_3 ? _matrix_b_4_T_10 : _GEN_6412; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 254:24 284:27]
  wire [255:0] _GEN_6432 = _T_3 ? _matrix_c_4_T_10 : _GEN_6417; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 254:24 285:27]
  wire [255:0] _GEN_6449 = _T_2 ? _GEN_6400 : _GEN_6422; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 254:24]
  wire [255:0] _GEN_6454 = _T_2 ? _GEN_6401 : _GEN_6427; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 254:24]
  wire [255:0] _GEN_6459 = _T_2 ? _GEN_6402 : _GEN_6432; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 254:24]
  wire [63:0] a_tile_v_108_1 = rf_a_tile_v_1_MPORT_108_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] a_tile_v_108_0 = rf_a_tile_v_0_MPORT_108_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_a_4_T_8 = {a_tile_v_108_1,a_tile_v_108_0,128'h0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 300:35]
  wire [63:0] matrix_b_4_tile_v_12_3 = rf_matrix_b_4_tile_v_3_MPORT_12_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_4_tile_v_12_2 = rf_matrix_b_4_tile_v_2_MPORT_12_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_4_tile_v_12_1 = rf_matrix_b_4_tile_v_1_MPORT_12_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_4_tile_v_12_0 = rf_matrix_b_4_tile_v_0_MPORT_12_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_b_4_T_12 = {matrix_b_4_tile_v_12_3,matrix_b_4_tile_v_12_2,matrix_b_4_tile_v_12_1,
    matrix_b_4_tile_v_12_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] matrix_c_4_tile_v_12_3 = rf_matrix_c_4_tile_v_3_MPORT_12_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_4_tile_v_12_2 = rf_matrix_c_4_tile_v_2_MPORT_12_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_4_tile_v_12_1 = rf_matrix_c_4_tile_v_1_MPORT_12_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_4_tile_v_12_0 = rf_matrix_c_4_tile_v_0_MPORT_12_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_c_4_T_12 = {matrix_c_4_tile_v_12_3,matrix_c_4_tile_v_12_2,matrix_c_4_tile_v_12_1,
    matrix_c_4_tile_v_12_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] a_tile_v_109_3 = rf_a_tile_v_3_MPORT_36_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] a_tile_v_109_2 = rf_a_tile_v_2_MPORT_36_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] a_tile_v_109_1 = rf_a_tile_v_1_MPORT_109_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] a_tile_v_109_0 = rf_a_tile_v_0_MPORT_109_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] a_109 = {a_tile_v_109_3,a_tile_v_109_2,a_tile_v_109_1,a_tile_v_109_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] matrix_b_4_tile_v_13_3 = rf_matrix_b_4_tile_v_3_MPORT_13_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_4_tile_v_13_2 = rf_matrix_b_4_tile_v_2_MPORT_13_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_4_tile_v_13_1 = rf_matrix_b_4_tile_v_1_MPORT_13_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_4_tile_v_13_0 = rf_matrix_b_4_tile_v_0_MPORT_13_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_b_4_T_13 = {matrix_b_4_tile_v_13_3,matrix_b_4_tile_v_13_2,matrix_b_4_tile_v_13_1,
    matrix_b_4_tile_v_13_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] matrix_c_4_tile_v_13_3 = rf_matrix_c_4_tile_v_3_MPORT_13_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_4_tile_v_13_2 = rf_matrix_c_4_tile_v_2_MPORT_13_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_4_tile_v_13_1 = rf_matrix_c_4_tile_v_1_MPORT_13_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_4_tile_v_13_0 = rf_matrix_c_4_tile_v_0_MPORT_13_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_c_4_T_13 = {matrix_c_4_tile_v_13_3,matrix_c_4_tile_v_13_2,matrix_c_4_tile_v_13_1,
    matrix_c_4_tile_v_13_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [255:0] _GEN_6579 = io_mixPc ? _matrix_a_4_T_8 : a_109; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 298:30 300:29 305:29]
  wire [255:0] _GEN_6584 = io_mixPc ? _matrix_b_4_T_12 : _matrix_b_4_T_13; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 298:30 301:29 306:29]
  wire [255:0] _GEN_6585 = io_mixPc ? _matrix_c_4_T_12 : _matrix_c_4_T_13; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 298:30 302:29 307:29]
  wire [63:0] a_tile_v_110_1 = rf_a_tile_v_1_MPORT_110_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] a_tile_v_110_0 = rf_a_tile_v_0_MPORT_110_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_a_4_T_9 = {a_tile_v_110_1,a_tile_v_110_0,128'h0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 313:35]
  wire [63:0] matrix_b_4_tile_v_14_3 = rf_matrix_b_4_tile_v_3_MPORT_14_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_4_tile_v_14_2 = rf_matrix_b_4_tile_v_2_MPORT_14_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_4_tile_v_14_1 = rf_matrix_b_4_tile_v_1_MPORT_14_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_4_tile_v_14_0 = rf_matrix_b_4_tile_v_0_MPORT_14_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_b_4_T_14 = {matrix_b_4_tile_v_14_3,matrix_b_4_tile_v_14_2,matrix_b_4_tile_v_14_1,
    matrix_b_4_tile_v_14_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] matrix_c_4_tile_v_14_3 = rf_matrix_c_4_tile_v_3_MPORT_14_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_4_tile_v_14_2 = rf_matrix_c_4_tile_v_2_MPORT_14_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_4_tile_v_14_1 = rf_matrix_c_4_tile_v_1_MPORT_14_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_4_tile_v_14_0 = rf_matrix_c_4_tile_v_0_MPORT_14_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_c_4_T_14 = {matrix_c_4_tile_v_14_3,matrix_c_4_tile_v_14_2,matrix_c_4_tile_v_14_1,
    matrix_c_4_tile_v_14_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] a_tile_v_111_3 = rf_a_tile_v_3_MPORT_37_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] a_tile_v_111_2 = rf_a_tile_v_2_MPORT_37_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] a_tile_v_111_1 = rf_a_tile_v_1_MPORT_111_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] a_tile_v_111_0 = rf_a_tile_v_0_MPORT_111_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] a_111 = {a_tile_v_111_3,a_tile_v_111_2,a_tile_v_111_1,a_tile_v_111_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] matrix_b_4_tile_v_15_3 = rf_matrix_b_4_tile_v_3_MPORT_15_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_4_tile_v_15_2 = rf_matrix_b_4_tile_v_2_MPORT_15_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_4_tile_v_15_1 = rf_matrix_b_4_tile_v_1_MPORT_15_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_4_tile_v_15_0 = rf_matrix_b_4_tile_v_0_MPORT_15_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_b_4_T_15 = {matrix_b_4_tile_v_15_3,matrix_b_4_tile_v_15_2,matrix_b_4_tile_v_15_1,
    matrix_b_4_tile_v_15_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] matrix_c_4_tile_v_15_3 = rf_matrix_c_4_tile_v_3_MPORT_15_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_4_tile_v_15_2 = rf_matrix_c_4_tile_v_2_MPORT_15_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_4_tile_v_15_1 = rf_matrix_c_4_tile_v_1_MPORT_15_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_4_tile_v_15_0 = rf_matrix_c_4_tile_v_0_MPORT_15_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_c_4_T_15 = {matrix_c_4_tile_v_15_3,matrix_c_4_tile_v_15_2,matrix_c_4_tile_v_15_1,
    matrix_c_4_tile_v_15_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [255:0] _GEN_6596 = io_mixPc ? _matrix_a_4_T_9 : a_111; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 311:30 313:29 318:29]
  wire [255:0] _GEN_6597 = io_mixPc ? _matrix_b_4_T_14 : _matrix_b_4_T_15; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 311:30 314:29 319:29]
  wire [255:0] _GEN_6598 = io_mixPc ? _matrix_c_4_T_14 : _matrix_c_4_T_15; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 311:30 315:29 320:29]
  wire [63:0] a_tile_v_112_1 = rf_a_tile_v_1_MPORT_112_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] a_tile_v_112_0 = rf_a_tile_v_0_MPORT_112_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_a_4_T_10 = {a_tile_v_112_1,a_tile_v_112_0,128'h0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 325:33]
  wire [63:0] matrix_b_4_tile_v_16_3 = rf_matrix_b_4_tile_v_3_MPORT_16_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_4_tile_v_16_2 = rf_matrix_b_4_tile_v_2_MPORT_16_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_4_tile_v_16_1 = rf_matrix_b_4_tile_v_1_MPORT_16_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_4_tile_v_16_0 = rf_matrix_b_4_tile_v_0_MPORT_16_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_b_4_T_16 = {matrix_b_4_tile_v_16_3,matrix_b_4_tile_v_16_2,matrix_b_4_tile_v_16_1,
    matrix_b_4_tile_v_16_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] matrix_c_4_tile_v_16_3 = rf_matrix_c_4_tile_v_3_MPORT_16_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_4_tile_v_16_2 = rf_matrix_c_4_tile_v_2_MPORT_16_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_4_tile_v_16_1 = rf_matrix_c_4_tile_v_1_MPORT_16_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_4_tile_v_16_0 = rf_matrix_c_4_tile_v_0_MPORT_16_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_c_4_T_16 = {matrix_c_4_tile_v_16_3,matrix_c_4_tile_v_16_2,matrix_c_4_tile_v_16_1,
    matrix_c_4_tile_v_16_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] a_tile_v_113_1 = rf_a_tile_v_1_MPORT_113_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] a_tile_v_113_0 = rf_a_tile_v_0_MPORT_113_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_a_4_T_11 = {a_tile_v_113_1,a_tile_v_113_0,128'h0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 331:33]
  wire [63:0] matrix_b_4_tile_v_17_3 = rf_matrix_b_4_tile_v_3_MPORT_17_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_4_tile_v_17_2 = rf_matrix_b_4_tile_v_2_MPORT_17_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_4_tile_v_17_1 = rf_matrix_b_4_tile_v_1_MPORT_17_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_4_tile_v_17_0 = rf_matrix_b_4_tile_v_0_MPORT_17_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_b_4_T_17 = {matrix_b_4_tile_v_17_3,matrix_b_4_tile_v_17_2,matrix_b_4_tile_v_17_1,
    matrix_b_4_tile_v_17_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] matrix_c_4_tile_v_17_3 = rf_matrix_c_4_tile_v_3_MPORT_17_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_4_tile_v_17_2 = rf_matrix_c_4_tile_v_2_MPORT_17_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_4_tile_v_17_1 = rf_matrix_c_4_tile_v_1_MPORT_17_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_4_tile_v_17_0 = rf_matrix_c_4_tile_v_0_MPORT_17_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_c_4_T_17 = {matrix_c_4_tile_v_17_3,matrix_c_4_tile_v_17_2,matrix_c_4_tile_v_17_1,
    matrix_c_4_tile_v_17_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [255:0] _GEN_6603 = _T_4 ? _matrix_a_4_T_11 : matrix_a_4; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 159:21 296:24 331:27]
  wire [255:0] _GEN_6608 = _T_4 ? _matrix_b_4_T_17 : matrix_b_4; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 160:21 296:24 332:27]
  wire [255:0] _GEN_6613 = _T_4 ? _matrix_c_4_T_17 : matrix_c_4; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 161:21 296:24 333:27]
  wire [255:0] _GEN_6618 = _T_3 ? _matrix_a_4_T_10 : _GEN_6603; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 296:24 325:27]
  wire [255:0] _GEN_6623 = _T_3 ? _matrix_b_4_T_16 : _GEN_6608; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 296:24 326:27]
  wire [255:0] _GEN_6628 = _T_3 ? _matrix_c_4_T_16 : _GEN_6613; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 296:24 327:27]
  wire [255:0] _GEN_6645 = _T_2 ? _GEN_6596 : _GEN_6618; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 296:24]
  wire [255:0] _GEN_6650 = _T_2 ? _GEN_6597 : _GEN_6623; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 296:24]
  wire [255:0] _GEN_6655 = _T_2 ? _GEN_6598 : _GEN_6628; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 296:24]
  wire [255:0] _GEN_6698 = _T_1 ? _GEN_6579 : _GEN_6645; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 296:24]
  wire [255:0] _GEN_6703 = _T_1 ? _GEN_6584 : _GEN_6650; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 296:24]
  wire [255:0] _GEN_6708 = _T_1 ? _GEN_6585 : _GEN_6655; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 296:24]
  wire [63:0] a_tile_v_114_1 = rf_a_tile_v_1_MPORT_114_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] a_tile_v_114_0 = rf_a_tile_v_0_MPORT_114_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_a_4_T_12 = {a_tile_v_114_1,a_tile_v_114_0,128'h0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 342:35]
  wire [63:0] matrix_b_4_tile_v_18_3 = rf_matrix_b_4_tile_v_3_MPORT_18_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_4_tile_v_18_2 = rf_matrix_b_4_tile_v_2_MPORT_18_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_4_tile_v_18_1 = rf_matrix_b_4_tile_v_1_MPORT_18_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_4_tile_v_18_0 = rf_matrix_b_4_tile_v_0_MPORT_18_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_b_4_T_18 = {matrix_b_4_tile_v_18_3,matrix_b_4_tile_v_18_2,matrix_b_4_tile_v_18_1,
    matrix_b_4_tile_v_18_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] matrix_c_4_tile_v_18_3 = rf_matrix_c_4_tile_v_3_MPORT_18_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_4_tile_v_18_2 = rf_matrix_c_4_tile_v_2_MPORT_18_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_4_tile_v_18_1 = rf_matrix_c_4_tile_v_1_MPORT_18_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_4_tile_v_18_0 = rf_matrix_c_4_tile_v_0_MPORT_18_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_c_4_T_18 = {matrix_c_4_tile_v_18_3,matrix_c_4_tile_v_18_2,matrix_c_4_tile_v_18_1,
    matrix_c_4_tile_v_18_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] a_tile_v_115_3 = rf_a_tile_v_3_MPORT_38_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] a_tile_v_115_2 = rf_a_tile_v_2_MPORT_38_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] a_tile_v_115_1 = rf_a_tile_v_1_MPORT_115_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] a_tile_v_115_0 = rf_a_tile_v_0_MPORT_115_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] a_115 = {a_tile_v_115_3,a_tile_v_115_2,a_tile_v_115_1,a_tile_v_115_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] matrix_b_4_tile_v_19_3 = rf_matrix_b_4_tile_v_3_MPORT_19_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_4_tile_v_19_2 = rf_matrix_b_4_tile_v_2_MPORT_19_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_4_tile_v_19_1 = rf_matrix_b_4_tile_v_1_MPORT_19_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_4_tile_v_19_0 = rf_matrix_b_4_tile_v_0_MPORT_19_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_b_4_T_19 = {matrix_b_4_tile_v_19_3,matrix_b_4_tile_v_19_2,matrix_b_4_tile_v_19_1,
    matrix_b_4_tile_v_19_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] matrix_c_4_tile_v_19_3 = rf_matrix_c_4_tile_v_3_MPORT_19_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_4_tile_v_19_2 = rf_matrix_c_4_tile_v_2_MPORT_19_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_4_tile_v_19_1 = rf_matrix_c_4_tile_v_1_MPORT_19_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_4_tile_v_19_0 = rf_matrix_c_4_tile_v_0_MPORT_19_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_c_4_T_19 = {matrix_c_4_tile_v_19_3,matrix_c_4_tile_v_19_2,matrix_c_4_tile_v_19_1,
    matrix_c_4_tile_v_19_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [255:0] _GEN_6775 = io_mixPc ? _matrix_a_4_T_12 : a_115; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 340:30 342:29 347:29]
  wire [255:0] _GEN_6780 = io_mixPc ? _matrix_b_4_T_18 : _matrix_b_4_T_19; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 340:30 343:29 348:29]
  wire [255:0] _GEN_6781 = io_mixPc ? _matrix_c_4_T_18 : _matrix_c_4_T_19; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 340:30 344:29 349:29]
  wire [63:0] a_tile_v_116_1 = rf_a_tile_v_1_MPORT_116_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] a_tile_v_116_0 = rf_a_tile_v_0_MPORT_116_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_a_4_T_13 = {a_tile_v_116_1,a_tile_v_116_0,128'h0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 355:35]
  wire [63:0] matrix_b_4_tile_v_20_3 = rf_matrix_b_4_tile_v_3_MPORT_20_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_4_tile_v_20_2 = rf_matrix_b_4_tile_v_2_MPORT_20_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_4_tile_v_20_1 = rf_matrix_b_4_tile_v_1_MPORT_20_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_4_tile_v_20_0 = rf_matrix_b_4_tile_v_0_MPORT_20_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_b_4_T_20 = {matrix_b_4_tile_v_20_3,matrix_b_4_tile_v_20_2,matrix_b_4_tile_v_20_1,
    matrix_b_4_tile_v_20_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] matrix_c_4_tile_v_20_3 = rf_matrix_c_4_tile_v_3_MPORT_20_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_4_tile_v_20_2 = rf_matrix_c_4_tile_v_2_MPORT_20_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_4_tile_v_20_1 = rf_matrix_c_4_tile_v_1_MPORT_20_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_4_tile_v_20_0 = rf_matrix_c_4_tile_v_0_MPORT_20_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_c_4_T_20 = {matrix_c_4_tile_v_20_3,matrix_c_4_tile_v_20_2,matrix_c_4_tile_v_20_1,
    matrix_c_4_tile_v_20_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] a_tile_v_117_3 = rf_a_tile_v_3_MPORT_39_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] a_tile_v_117_2 = rf_a_tile_v_2_MPORT_39_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] a_tile_v_117_1 = rf_a_tile_v_1_MPORT_117_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] a_tile_v_117_0 = rf_a_tile_v_0_MPORT_117_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] a_117 = {a_tile_v_117_3,a_tile_v_117_2,a_tile_v_117_1,a_tile_v_117_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] matrix_b_4_tile_v_21_3 = rf_matrix_b_4_tile_v_3_MPORT_21_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_4_tile_v_21_2 = rf_matrix_b_4_tile_v_2_MPORT_21_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_4_tile_v_21_1 = rf_matrix_b_4_tile_v_1_MPORT_21_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_4_tile_v_21_0 = rf_matrix_b_4_tile_v_0_MPORT_21_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_b_4_T_21 = {matrix_b_4_tile_v_21_3,matrix_b_4_tile_v_21_2,matrix_b_4_tile_v_21_1,
    matrix_b_4_tile_v_21_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] matrix_c_4_tile_v_21_3 = rf_matrix_c_4_tile_v_3_MPORT_21_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_4_tile_v_21_2 = rf_matrix_c_4_tile_v_2_MPORT_21_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_4_tile_v_21_1 = rf_matrix_c_4_tile_v_1_MPORT_21_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_4_tile_v_21_0 = rf_matrix_c_4_tile_v_0_MPORT_21_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_c_4_T_21 = {matrix_c_4_tile_v_21_3,matrix_c_4_tile_v_21_2,matrix_c_4_tile_v_21_1,
    matrix_c_4_tile_v_21_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [255:0] _GEN_6792 = io_mixPc ? _matrix_a_4_T_13 : a_117; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 353:30 355:29 360:29]
  wire [255:0] _GEN_6793 = io_mixPc ? _matrix_b_4_T_20 : _matrix_b_4_T_21; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 353:30 356:29 361:29]
  wire [255:0] _GEN_6794 = io_mixPc ? _matrix_c_4_T_20 : _matrix_c_4_T_21; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 353:30 357:29 362:29]
  wire [63:0] a_tile_v_118_1 = rf_a_tile_v_1_MPORT_118_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] a_tile_v_118_0 = rf_a_tile_v_0_MPORT_118_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_a_4_T_14 = {a_tile_v_118_1,a_tile_v_118_0,128'h0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 367:33]
  wire [63:0] matrix_b_4_tile_v_22_3 = rf_matrix_b_4_tile_v_3_MPORT_22_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_4_tile_v_22_2 = rf_matrix_b_4_tile_v_2_MPORT_22_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_4_tile_v_22_1 = rf_matrix_b_4_tile_v_1_MPORT_22_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_4_tile_v_22_0 = rf_matrix_b_4_tile_v_0_MPORT_22_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_b_4_T_22 = {matrix_b_4_tile_v_22_3,matrix_b_4_tile_v_22_2,matrix_b_4_tile_v_22_1,
    matrix_b_4_tile_v_22_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] matrix_c_4_tile_v_22_3 = rf_matrix_c_4_tile_v_3_MPORT_22_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_4_tile_v_22_2 = rf_matrix_c_4_tile_v_2_MPORT_22_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_4_tile_v_22_1 = rf_matrix_c_4_tile_v_1_MPORT_22_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_4_tile_v_22_0 = rf_matrix_c_4_tile_v_0_MPORT_22_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_c_4_T_22 = {matrix_c_4_tile_v_22_3,matrix_c_4_tile_v_22_2,matrix_c_4_tile_v_22_1,
    matrix_c_4_tile_v_22_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] a_tile_v_119_1 = rf_a_tile_v_1_MPORT_119_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] a_tile_v_119_0 = rf_a_tile_v_0_MPORT_119_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_a_4_T_15 = {a_tile_v_119_1,a_tile_v_119_0,128'h0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 373:33]
  wire [63:0] matrix_b_4_tile_v_23_3 = rf_matrix_b_4_tile_v_3_MPORT_23_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_4_tile_v_23_2 = rf_matrix_b_4_tile_v_2_MPORT_23_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_4_tile_v_23_1 = rf_matrix_b_4_tile_v_1_MPORT_23_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_4_tile_v_23_0 = rf_matrix_b_4_tile_v_0_MPORT_23_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_b_4_T_23 = {matrix_b_4_tile_v_23_3,matrix_b_4_tile_v_23_2,matrix_b_4_tile_v_23_1,
    matrix_b_4_tile_v_23_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] matrix_c_4_tile_v_23_3 = rf_matrix_c_4_tile_v_3_MPORT_23_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_4_tile_v_23_2 = rf_matrix_c_4_tile_v_2_MPORT_23_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_4_tile_v_23_1 = rf_matrix_c_4_tile_v_1_MPORT_23_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_4_tile_v_23_0 = rf_matrix_c_4_tile_v_0_MPORT_23_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_c_4_T_23 = {matrix_c_4_tile_v_23_3,matrix_c_4_tile_v_23_2,matrix_c_4_tile_v_23_1,
    matrix_c_4_tile_v_23_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [255:0] _GEN_6799 = _T_4 ? _matrix_a_4_T_15 : matrix_a_4; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 159:21 338:24 373:27]
  wire [255:0] _GEN_6804 = _T_4 ? _matrix_b_4_T_23 : matrix_b_4; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 160:21 338:24 374:27]
  wire [255:0] _GEN_6809 = _T_4 ? _matrix_c_4_T_23 : matrix_c_4; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 161:21 338:24 375:27]
  wire [255:0] _GEN_6814 = _T_3 ? _matrix_a_4_T_14 : _GEN_6799; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 338:24 367:27]
  wire [255:0] _GEN_6819 = _T_3 ? _matrix_b_4_T_22 : _GEN_6804; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 338:24 368:27]
  wire [255:0] _GEN_6824 = _T_3 ? _matrix_c_4_T_22 : _GEN_6809; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 338:24 369:27]
  wire [255:0] _GEN_6841 = _T_2 ? _GEN_6792 : _GEN_6814; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 338:24]
  wire [255:0] _GEN_6846 = _T_2 ? _GEN_6793 : _GEN_6819; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 338:24]
  wire [255:0] _GEN_6851 = _T_2 ? _GEN_6794 : _GEN_6824; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 338:24]
  wire [255:0] _GEN_6894 = _T_1 ? _GEN_6775 : _GEN_6841; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 338:24]
  wire [255:0] _GEN_6899 = _T_1 ? _GEN_6780 : _GEN_6846; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 338:24]
  wire [255:0] _GEN_6904 = _T_1 ? _GEN_6781 : _GEN_6851; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 338:24]
  wire [255:0] _GEN_6973 = 2'h3 == set ? _GEN_6894 : matrix_a_4; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 210:18 159:21]
  wire [255:0] _GEN_6978 = 2'h3 == set ? _GEN_6899 : matrix_b_4; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 210:18 160:21]
  wire [255:0] _GEN_6983 = 2'h3 == set ? _GEN_6904 : matrix_c_4; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 210:18 161:21]
  wire [63:0] a_tile_v_120_1 = rf_a_tile_v_1_MPORT_120_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] a_tile_v_120_0 = rf_a_tile_v_0_MPORT_120_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_a_5_T = {a_tile_v_120_1,a_tile_v_120_0,128'h0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 216:35]
  wire [63:0] matrix_b_5_tile_v__3 = rf_matrix_b_5_tile_v_3_MPORT_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_5_tile_v__2 = rf_matrix_b_5_tile_v_2_MPORT_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_5_tile_v__1 = rf_matrix_b_5_tile_v_1_MPORT_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_5_tile_v__0 = rf_matrix_b_5_tile_v_0_MPORT_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_b_5_T = {matrix_b_5_tile_v__3,matrix_b_5_tile_v__2,matrix_b_5_tile_v__1,matrix_b_5_tile_v__0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] matrix_c_5_tile_v__3 = rf_matrix_c_5_tile_v_3_MPORT_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_5_tile_v__2 = rf_matrix_c_5_tile_v_2_MPORT_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_5_tile_v__1 = rf_matrix_c_5_tile_v_1_MPORT_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_5_tile_v__0 = rf_matrix_c_5_tile_v_0_MPORT_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_c_5_T = {matrix_c_5_tile_v__3,matrix_c_5_tile_v__2,matrix_c_5_tile_v__1,matrix_c_5_tile_v__0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] a_tile_v_121_3 = rf_a_tile_v_3_MPORT_40_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] a_tile_v_121_2 = rf_a_tile_v_2_MPORT_40_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] a_tile_v_121_1 = rf_a_tile_v_1_MPORT_121_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] a_tile_v_121_0 = rf_a_tile_v_0_MPORT_121_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] a_121 = {a_tile_v_121_3,a_tile_v_121_2,a_tile_v_121_1,a_tile_v_121_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] matrix_b_5_tile_v_1_3 = rf_matrix_b_5_tile_v_3_MPORT_1_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_5_tile_v_1_2 = rf_matrix_b_5_tile_v_2_MPORT_1_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_5_tile_v_1_1 = rf_matrix_b_5_tile_v_1_MPORT_1_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_5_tile_v_1_0 = rf_matrix_b_5_tile_v_0_MPORT_1_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_b_5_T_1 = {matrix_b_5_tile_v_1_3,matrix_b_5_tile_v_1_2,matrix_b_5_tile_v_1_1,
    matrix_b_5_tile_v_1_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] matrix_c_5_tile_v_1_3 = rf_matrix_c_5_tile_v_3_MPORT_1_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_5_tile_v_1_2 = rf_matrix_c_5_tile_v_2_MPORT_1_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_5_tile_v_1_1 = rf_matrix_c_5_tile_v_1_MPORT_1_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_5_tile_v_1_0 = rf_matrix_c_5_tile_v_0_MPORT_1_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_c_5_T_1 = {matrix_c_5_tile_v_1_3,matrix_c_5_tile_v_1_2,matrix_c_5_tile_v_1_1,
    matrix_c_5_tile_v_1_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] a_tile_v_122_1 = rf_a_tile_v_1_MPORT_122_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] a_tile_v_122_0 = rf_a_tile_v_0_MPORT_122_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_a_5_T_1 = {a_tile_v_122_1,a_tile_v_122_0,128'h0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 229:35]
  wire [63:0] matrix_b_5_tile_v_2_3 = rf_matrix_b_5_tile_v_3_MPORT_2_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_5_tile_v_2_2 = rf_matrix_b_5_tile_v_2_MPORT_2_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_5_tile_v_2_1 = rf_matrix_b_5_tile_v_1_MPORT_2_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_5_tile_v_2_0 = rf_matrix_b_5_tile_v_0_MPORT_2_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_b_5_T_2 = {matrix_b_5_tile_v_2_3,matrix_b_5_tile_v_2_2,matrix_b_5_tile_v_2_1,
    matrix_b_5_tile_v_2_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] matrix_c_5_tile_v_2_3 = rf_matrix_c_5_tile_v_3_MPORT_2_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_5_tile_v_2_2 = rf_matrix_c_5_tile_v_2_MPORT_2_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_5_tile_v_2_1 = rf_matrix_c_5_tile_v_1_MPORT_2_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_5_tile_v_2_0 = rf_matrix_c_5_tile_v_0_MPORT_2_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_c_5_T_2 = {matrix_c_5_tile_v_2_3,matrix_c_5_tile_v_2_2,matrix_c_5_tile_v_2_1,
    matrix_c_5_tile_v_2_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] a_tile_v_123_3 = rf_a_tile_v_3_MPORT_41_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] a_tile_v_123_2 = rf_a_tile_v_2_MPORT_41_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] a_tile_v_123_1 = rf_a_tile_v_1_MPORT_123_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] a_tile_v_123_0 = rf_a_tile_v_0_MPORT_123_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] a_123 = {a_tile_v_123_3,a_tile_v_123_2,a_tile_v_123_1,a_tile_v_123_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] matrix_b_5_tile_v_3_3 = rf_matrix_b_5_tile_v_3_MPORT_3_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_5_tile_v_3_2 = rf_matrix_b_5_tile_v_2_MPORT_3_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_5_tile_v_3_1 = rf_matrix_b_5_tile_v_1_MPORT_3_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_5_tile_v_3_0 = rf_matrix_b_5_tile_v_0_MPORT_3_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_b_5_T_3 = {matrix_b_5_tile_v_3_3,matrix_b_5_tile_v_3_2,matrix_b_5_tile_v_3_1,
    matrix_b_5_tile_v_3_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] matrix_c_5_tile_v_3_3 = rf_matrix_c_5_tile_v_3_MPORT_3_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_5_tile_v_3_2 = rf_matrix_c_5_tile_v_2_MPORT_3_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_5_tile_v_3_1 = rf_matrix_c_5_tile_v_1_MPORT_3_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_5_tile_v_3_0 = rf_matrix_c_5_tile_v_0_MPORT_3_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_c_5_T_3 = {matrix_c_5_tile_v_3_3,matrix_c_5_tile_v_3_2,matrix_c_5_tile_v_3_1,
    matrix_c_5_tile_v_3_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [255:0] _GEN_7760 = io_mixPc ? _matrix_a_5_T_1 : a_123; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 227:30 229:29 234:29]
  wire [255:0] _GEN_7761 = io_mixPc ? _matrix_b_5_T_2 : _matrix_b_5_T_3; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 227:30 230:29 235:29]
  wire [255:0] _GEN_7766 = io_mixPc ? _matrix_c_5_T_2 : _matrix_c_5_T_3; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 227:30 231:29 236:29]
  wire [63:0] a_tile_v_124_1 = rf_a_tile_v_1_MPORT_124_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] a_tile_v_124_0 = rf_a_tile_v_0_MPORT_124_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_a_5_T_2 = {a_tile_v_124_1,a_tile_v_124_0,128'h0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 241:33]
  wire [63:0] matrix_b_5_tile_v_4_3 = rf_matrix_b_5_tile_v_3_MPORT_4_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_5_tile_v_4_2 = rf_matrix_b_5_tile_v_2_MPORT_4_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_5_tile_v_4_1 = rf_matrix_b_5_tile_v_1_MPORT_4_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_5_tile_v_4_0 = rf_matrix_b_5_tile_v_0_MPORT_4_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_b_5_T_4 = {matrix_b_5_tile_v_4_3,matrix_b_5_tile_v_4_2,matrix_b_5_tile_v_4_1,
    matrix_b_5_tile_v_4_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] matrix_c_5_tile_v_4_3 = rf_matrix_c_5_tile_v_3_MPORT_4_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_5_tile_v_4_2 = rf_matrix_c_5_tile_v_2_MPORT_4_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_5_tile_v_4_1 = rf_matrix_c_5_tile_v_1_MPORT_4_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_5_tile_v_4_0 = rf_matrix_c_5_tile_v_0_MPORT_4_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_c_5_T_4 = {matrix_c_5_tile_v_4_3,matrix_c_5_tile_v_4_2,matrix_c_5_tile_v_4_1,
    matrix_c_5_tile_v_4_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] a_tile_v_125_1 = rf_a_tile_v_1_MPORT_125_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] a_tile_v_125_0 = rf_a_tile_v_0_MPORT_125_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_a_5_T_3 = {a_tile_v_125_1,a_tile_v_125_0,128'h0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 247:33]
  wire [63:0] matrix_b_5_tile_v_5_3 = rf_matrix_b_5_tile_v_3_MPORT_5_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_5_tile_v_5_2 = rf_matrix_b_5_tile_v_2_MPORT_5_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_5_tile_v_5_1 = rf_matrix_b_5_tile_v_1_MPORT_5_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_5_tile_v_5_0 = rf_matrix_b_5_tile_v_0_MPORT_5_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_b_5_T_5 = {matrix_b_5_tile_v_5_3,matrix_b_5_tile_v_5_2,matrix_b_5_tile_v_5_1,
    matrix_b_5_tile_v_5_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] matrix_c_5_tile_v_5_3 = rf_matrix_c_5_tile_v_3_MPORT_5_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_5_tile_v_5_2 = rf_matrix_c_5_tile_v_2_MPORT_5_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_5_tile_v_5_1 = rf_matrix_c_5_tile_v_1_MPORT_5_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_5_tile_v_5_0 = rf_matrix_c_5_tile_v_0_MPORT_5_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_c_5_T_5 = {matrix_c_5_tile_v_5_3,matrix_c_5_tile_v_5_2,matrix_c_5_tile_v_5_1,
    matrix_c_5_tile_v_5_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [255:0] _GEN_7775 = 2'h3 == step ? _matrix_a_5_T_3 : matrix_a_5; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 159:21 212:23 247:27]
  wire [255:0] _GEN_7780 = 2'h3 == step ? _matrix_b_5_T_5 : matrix_b_5; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 160:21 212:23 248:27]
  wire [255:0] _GEN_7785 = 2'h3 == step ? _matrix_c_5_T_5 : matrix_c_5; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 161:21 212:23 249:27]
  wire [255:0] _GEN_7790 = 2'h2 == step ? _matrix_a_5_T_2 : _GEN_7775; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 212:23 241:27]
  wire [255:0] _GEN_7795 = 2'h2 == step ? _matrix_b_5_T_4 : _GEN_7780; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 212:23 242:27]
  wire [255:0] _GEN_7800 = 2'h2 == step ? _matrix_c_5_T_4 : _GEN_7785; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 212:23 243:27]
  wire [63:0] a_tile_v_126_1 = rf_a_tile_v_1_MPORT_126_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] a_tile_v_126_0 = rf_a_tile_v_0_MPORT_126_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_a_5_T_4 = {a_tile_v_126_1,a_tile_v_126_0,128'h0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 258:35]
  wire [63:0] matrix_b_5_tile_v_6_3 = rf_matrix_b_5_tile_v_3_MPORT_6_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_5_tile_v_6_2 = rf_matrix_b_5_tile_v_2_MPORT_6_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_5_tile_v_6_1 = rf_matrix_b_5_tile_v_1_MPORT_6_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_5_tile_v_6_0 = rf_matrix_b_5_tile_v_0_MPORT_6_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_b_5_T_6 = {matrix_b_5_tile_v_6_3,matrix_b_5_tile_v_6_2,matrix_b_5_tile_v_6_1,
    matrix_b_5_tile_v_6_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] matrix_c_5_tile_v_6_3 = rf_matrix_c_5_tile_v_3_MPORT_6_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_5_tile_v_6_2 = rf_matrix_c_5_tile_v_2_MPORT_6_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_5_tile_v_6_1 = rf_matrix_c_5_tile_v_1_MPORT_6_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_5_tile_v_6_0 = rf_matrix_c_5_tile_v_0_MPORT_6_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_c_5_T_6 = {matrix_c_5_tile_v_6_3,matrix_c_5_tile_v_6_2,matrix_c_5_tile_v_6_1,
    matrix_c_5_tile_v_6_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] a_tile_v_127_3 = rf_a_tile_v_3_MPORT_42_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] a_tile_v_127_2 = rf_a_tile_v_2_MPORT_42_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] a_tile_v_127_1 = rf_a_tile_v_1_MPORT_127_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] a_tile_v_127_0 = rf_a_tile_v_0_MPORT_127_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] a_127 = {a_tile_v_127_3,a_tile_v_127_2,a_tile_v_127_1,a_tile_v_127_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] matrix_b_5_tile_v_7_3 = rf_matrix_b_5_tile_v_3_MPORT_7_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_5_tile_v_7_2 = rf_matrix_b_5_tile_v_2_MPORT_7_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_5_tile_v_7_1 = rf_matrix_b_5_tile_v_1_MPORT_7_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_5_tile_v_7_0 = rf_matrix_b_5_tile_v_0_MPORT_7_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_b_5_T_7 = {matrix_b_5_tile_v_7_3,matrix_b_5_tile_v_7_2,matrix_b_5_tile_v_7_1,
    matrix_b_5_tile_v_7_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] matrix_c_5_tile_v_7_3 = rf_matrix_c_5_tile_v_3_MPORT_7_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_5_tile_v_7_2 = rf_matrix_c_5_tile_v_2_MPORT_7_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_5_tile_v_7_1 = rf_matrix_c_5_tile_v_1_MPORT_7_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_5_tile_v_7_0 = rf_matrix_c_5_tile_v_0_MPORT_7_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_c_5_T_7 = {matrix_c_5_tile_v_7_3,matrix_c_5_tile_v_7_2,matrix_c_5_tile_v_7_1,
    matrix_c_5_tile_v_7_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [255:0] _GEN_7947 = io_mixPc ? _matrix_a_5_T_4 : a_127; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 256:30 258:29 263:29]
  wire [255:0] _GEN_7948 = io_mixPc ? _matrix_b_5_T_6 : _matrix_b_5_T_7; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 256:30 259:29 264:29]
  wire [255:0] _GEN_7949 = io_mixPc ? _matrix_c_5_T_6 : _matrix_c_5_T_7; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 256:30 260:29 265:29]
  wire [63:0] a_tile_v_128_1 = rf_a_tile_v_1_MPORT_128_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] a_tile_v_128_0 = rf_a_tile_v_0_MPORT_128_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_a_5_T_5 = {a_tile_v_128_1,a_tile_v_128_0,128'h0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 271:35]
  wire [63:0] matrix_b_5_tile_v_8_3 = rf_matrix_b_5_tile_v_3_MPORT_8_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_5_tile_v_8_2 = rf_matrix_b_5_tile_v_2_MPORT_8_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_5_tile_v_8_1 = rf_matrix_b_5_tile_v_1_MPORT_8_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_5_tile_v_8_0 = rf_matrix_b_5_tile_v_0_MPORT_8_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_b_5_T_8 = {matrix_b_5_tile_v_8_3,matrix_b_5_tile_v_8_2,matrix_b_5_tile_v_8_1,
    matrix_b_5_tile_v_8_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] matrix_c_5_tile_v_8_3 = rf_matrix_c_5_tile_v_3_MPORT_8_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_5_tile_v_8_2 = rf_matrix_c_5_tile_v_2_MPORT_8_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_5_tile_v_8_1 = rf_matrix_c_5_tile_v_1_MPORT_8_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_5_tile_v_8_0 = rf_matrix_c_5_tile_v_0_MPORT_8_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_c_5_T_8 = {matrix_c_5_tile_v_8_3,matrix_c_5_tile_v_8_2,matrix_c_5_tile_v_8_1,
    matrix_c_5_tile_v_8_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] a_tile_v_129_3 = rf_a_tile_v_3_MPORT_43_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] a_tile_v_129_2 = rf_a_tile_v_2_MPORT_43_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] a_tile_v_129_1 = rf_a_tile_v_1_MPORT_129_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] a_tile_v_129_0 = rf_a_tile_v_0_MPORT_129_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] a_129 = {a_tile_v_129_3,a_tile_v_129_2,a_tile_v_129_1,a_tile_v_129_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] matrix_b_5_tile_v_9_3 = rf_matrix_b_5_tile_v_3_MPORT_9_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_5_tile_v_9_2 = rf_matrix_b_5_tile_v_2_MPORT_9_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_5_tile_v_9_1 = rf_matrix_b_5_tile_v_1_MPORT_9_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_5_tile_v_9_0 = rf_matrix_b_5_tile_v_0_MPORT_9_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_b_5_T_9 = {matrix_b_5_tile_v_9_3,matrix_b_5_tile_v_9_2,matrix_b_5_tile_v_9_1,
    matrix_b_5_tile_v_9_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] matrix_c_5_tile_v_9_3 = rf_matrix_c_5_tile_v_3_MPORT_9_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_5_tile_v_9_2 = rf_matrix_c_5_tile_v_2_MPORT_9_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_5_tile_v_9_1 = rf_matrix_c_5_tile_v_1_MPORT_9_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_5_tile_v_9_0 = rf_matrix_c_5_tile_v_0_MPORT_9_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_c_5_T_9 = {matrix_c_5_tile_v_9_3,matrix_c_5_tile_v_9_2,matrix_c_5_tile_v_9_1,
    matrix_c_5_tile_v_9_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [255:0] _GEN_7956 = io_mixPc ? _matrix_a_5_T_5 : a_129; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 269:30 271:29 276:29]
  wire [255:0] _GEN_7957 = io_mixPc ? _matrix_b_5_T_8 : _matrix_b_5_T_9; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 269:30 272:29 277:29]
  wire [255:0] _GEN_7958 = io_mixPc ? _matrix_c_5_T_8 : _matrix_c_5_T_9; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 269:30 273:29 278:29]
  wire [63:0] a_tile_v_130_1 = rf_a_tile_v_1_MPORT_130_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] a_tile_v_130_0 = rf_a_tile_v_0_MPORT_130_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_a_5_T_6 = {a_tile_v_130_1,a_tile_v_130_0,128'h0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 283:33]
  wire [63:0] matrix_b_5_tile_v_10_3 = rf_matrix_b_5_tile_v_3_MPORT_10_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_5_tile_v_10_2 = rf_matrix_b_5_tile_v_2_MPORT_10_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_5_tile_v_10_1 = rf_matrix_b_5_tile_v_1_MPORT_10_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_5_tile_v_10_0 = rf_matrix_b_5_tile_v_0_MPORT_10_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_b_5_T_10 = {matrix_b_5_tile_v_10_3,matrix_b_5_tile_v_10_2,matrix_b_5_tile_v_10_1,
    matrix_b_5_tile_v_10_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] matrix_c_5_tile_v_10_3 = rf_matrix_c_5_tile_v_3_MPORT_10_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_5_tile_v_10_2 = rf_matrix_c_5_tile_v_2_MPORT_10_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_5_tile_v_10_1 = rf_matrix_c_5_tile_v_1_MPORT_10_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_5_tile_v_10_0 = rf_matrix_c_5_tile_v_0_MPORT_10_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_c_5_T_10 = {matrix_c_5_tile_v_10_3,matrix_c_5_tile_v_10_2,matrix_c_5_tile_v_10_1,
    matrix_c_5_tile_v_10_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] a_tile_v_131_1 = rf_a_tile_v_1_MPORT_131_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] a_tile_v_131_0 = rf_a_tile_v_0_MPORT_131_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_a_5_T_7 = {a_tile_v_131_1,a_tile_v_131_0,128'h0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 289:33]
  wire [63:0] matrix_b_5_tile_v_11_3 = rf_matrix_b_5_tile_v_3_MPORT_11_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_5_tile_v_11_2 = rf_matrix_b_5_tile_v_2_MPORT_11_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_5_tile_v_11_1 = rf_matrix_b_5_tile_v_1_MPORT_11_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_5_tile_v_11_0 = rf_matrix_b_5_tile_v_0_MPORT_11_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_b_5_T_11 = {matrix_b_5_tile_v_11_3,matrix_b_5_tile_v_11_2,matrix_b_5_tile_v_11_1,
    matrix_b_5_tile_v_11_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] matrix_c_5_tile_v_11_3 = rf_matrix_c_5_tile_v_3_MPORT_11_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_5_tile_v_11_2 = rf_matrix_c_5_tile_v_2_MPORT_11_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_5_tile_v_11_1 = rf_matrix_c_5_tile_v_1_MPORT_11_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_5_tile_v_11_0 = rf_matrix_c_5_tile_v_0_MPORT_11_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_c_5_T_11 = {matrix_c_5_tile_v_11_3,matrix_c_5_tile_v_11_2,matrix_c_5_tile_v_11_1,
    matrix_c_5_tile_v_11_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [255:0] _GEN_7963 = _T_4 ? _matrix_a_5_T_7 : matrix_a_5; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 159:21 254:24 289:27]
  wire [255:0] _GEN_7968 = _T_4 ? _matrix_b_5_T_11 : matrix_b_5; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 160:21 254:24 290:27]
  wire [255:0] _GEN_7973 = _T_4 ? _matrix_c_5_T_11 : matrix_c_5; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 161:21 254:24 291:27]
  wire [255:0] _GEN_7978 = _T_3 ? _matrix_a_5_T_6 : _GEN_7963; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 254:24 283:27]
  wire [255:0] _GEN_7983 = _T_3 ? _matrix_b_5_T_10 : _GEN_7968; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 254:24 284:27]
  wire [255:0] _GEN_7988 = _T_3 ? _matrix_c_5_T_10 : _GEN_7973; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 254:24 285:27]
  wire [255:0] _GEN_8005 = _T_2 ? _GEN_7956 : _GEN_7978; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 254:24]
  wire [255:0] _GEN_8010 = _T_2 ? _GEN_7957 : _GEN_7983; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 254:24]
  wire [255:0] _GEN_8015 = _T_2 ? _GEN_7958 : _GEN_7988; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 254:24]
  wire [63:0] a_tile_v_132_1 = rf_a_tile_v_1_MPORT_132_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] a_tile_v_132_0 = rf_a_tile_v_0_MPORT_132_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_a_5_T_8 = {a_tile_v_132_1,a_tile_v_132_0,128'h0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 300:35]
  wire [63:0] matrix_b_5_tile_v_12_3 = rf_matrix_b_5_tile_v_3_MPORT_12_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_5_tile_v_12_2 = rf_matrix_b_5_tile_v_2_MPORT_12_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_5_tile_v_12_1 = rf_matrix_b_5_tile_v_1_MPORT_12_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_5_tile_v_12_0 = rf_matrix_b_5_tile_v_0_MPORT_12_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_b_5_T_12 = {matrix_b_5_tile_v_12_3,matrix_b_5_tile_v_12_2,matrix_b_5_tile_v_12_1,
    matrix_b_5_tile_v_12_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] matrix_c_5_tile_v_12_3 = rf_matrix_c_5_tile_v_3_MPORT_12_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_5_tile_v_12_2 = rf_matrix_c_5_tile_v_2_MPORT_12_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_5_tile_v_12_1 = rf_matrix_c_5_tile_v_1_MPORT_12_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_5_tile_v_12_0 = rf_matrix_c_5_tile_v_0_MPORT_12_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_c_5_T_12 = {matrix_c_5_tile_v_12_3,matrix_c_5_tile_v_12_2,matrix_c_5_tile_v_12_1,
    matrix_c_5_tile_v_12_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] a_tile_v_133_3 = rf_a_tile_v_3_MPORT_44_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] a_tile_v_133_2 = rf_a_tile_v_2_MPORT_44_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] a_tile_v_133_1 = rf_a_tile_v_1_MPORT_133_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] a_tile_v_133_0 = rf_a_tile_v_0_MPORT_133_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] a_133 = {a_tile_v_133_3,a_tile_v_133_2,a_tile_v_133_1,a_tile_v_133_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] matrix_b_5_tile_v_13_3 = rf_matrix_b_5_tile_v_3_MPORT_13_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_5_tile_v_13_2 = rf_matrix_b_5_tile_v_2_MPORT_13_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_5_tile_v_13_1 = rf_matrix_b_5_tile_v_1_MPORT_13_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_5_tile_v_13_0 = rf_matrix_b_5_tile_v_0_MPORT_13_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_b_5_T_13 = {matrix_b_5_tile_v_13_3,matrix_b_5_tile_v_13_2,matrix_b_5_tile_v_13_1,
    matrix_b_5_tile_v_13_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] matrix_c_5_tile_v_13_3 = rf_matrix_c_5_tile_v_3_MPORT_13_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_5_tile_v_13_2 = rf_matrix_c_5_tile_v_2_MPORT_13_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_5_tile_v_13_1 = rf_matrix_c_5_tile_v_1_MPORT_13_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_5_tile_v_13_0 = rf_matrix_c_5_tile_v_0_MPORT_13_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_c_5_T_13 = {matrix_c_5_tile_v_13_3,matrix_c_5_tile_v_13_2,matrix_c_5_tile_v_13_1,
    matrix_c_5_tile_v_13_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [255:0] _GEN_8135 = io_mixPc ? _matrix_a_5_T_8 : a_133; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 298:30 300:29 305:29]
  wire [255:0] _GEN_8136 = io_mixPc ? _matrix_b_5_T_12 : _matrix_b_5_T_13; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 298:30 301:29 306:29]
  wire [255:0] _GEN_8137 = io_mixPc ? _matrix_c_5_T_12 : _matrix_c_5_T_13; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 298:30 302:29 307:29]
  wire [63:0] a_tile_v_134_1 = rf_a_tile_v_1_MPORT_134_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] a_tile_v_134_0 = rf_a_tile_v_0_MPORT_134_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_a_5_T_9 = {a_tile_v_134_1,a_tile_v_134_0,128'h0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 313:35]
  wire [63:0] matrix_b_5_tile_v_14_3 = rf_matrix_b_5_tile_v_3_MPORT_14_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_5_tile_v_14_2 = rf_matrix_b_5_tile_v_2_MPORT_14_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_5_tile_v_14_1 = rf_matrix_b_5_tile_v_1_MPORT_14_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_5_tile_v_14_0 = rf_matrix_b_5_tile_v_0_MPORT_14_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_b_5_T_14 = {matrix_b_5_tile_v_14_3,matrix_b_5_tile_v_14_2,matrix_b_5_tile_v_14_1,
    matrix_b_5_tile_v_14_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] matrix_c_5_tile_v_14_3 = rf_matrix_c_5_tile_v_3_MPORT_14_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_5_tile_v_14_2 = rf_matrix_c_5_tile_v_2_MPORT_14_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_5_tile_v_14_1 = rf_matrix_c_5_tile_v_1_MPORT_14_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_5_tile_v_14_0 = rf_matrix_c_5_tile_v_0_MPORT_14_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_c_5_T_14 = {matrix_c_5_tile_v_14_3,matrix_c_5_tile_v_14_2,matrix_c_5_tile_v_14_1,
    matrix_c_5_tile_v_14_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] a_tile_v_135_3 = rf_a_tile_v_3_MPORT_45_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] a_tile_v_135_2 = rf_a_tile_v_2_MPORT_45_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] a_tile_v_135_1 = rf_a_tile_v_1_MPORT_135_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] a_tile_v_135_0 = rf_a_tile_v_0_MPORT_135_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] a_135 = {a_tile_v_135_3,a_tile_v_135_2,a_tile_v_135_1,a_tile_v_135_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] matrix_b_5_tile_v_15_3 = rf_matrix_b_5_tile_v_3_MPORT_15_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_5_tile_v_15_2 = rf_matrix_b_5_tile_v_2_MPORT_15_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_5_tile_v_15_1 = rf_matrix_b_5_tile_v_1_MPORT_15_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_5_tile_v_15_0 = rf_matrix_b_5_tile_v_0_MPORT_15_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_b_5_T_15 = {matrix_b_5_tile_v_15_3,matrix_b_5_tile_v_15_2,matrix_b_5_tile_v_15_1,
    matrix_b_5_tile_v_15_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] matrix_c_5_tile_v_15_3 = rf_matrix_c_5_tile_v_3_MPORT_15_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_5_tile_v_15_2 = rf_matrix_c_5_tile_v_2_MPORT_15_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_5_tile_v_15_1 = rf_matrix_c_5_tile_v_1_MPORT_15_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_5_tile_v_15_0 = rf_matrix_c_5_tile_v_0_MPORT_15_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_c_5_T_15 = {matrix_c_5_tile_v_15_3,matrix_c_5_tile_v_15_2,matrix_c_5_tile_v_15_1,
    matrix_c_5_tile_v_15_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [255:0] _GEN_8144 = io_mixPc ? _matrix_a_5_T_9 : a_135; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 311:30 313:29 318:29]
  wire [255:0] _GEN_8145 = io_mixPc ? _matrix_b_5_T_14 : _matrix_b_5_T_15; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 311:30 314:29 319:29]
  wire [255:0] _GEN_8146 = io_mixPc ? _matrix_c_5_T_14 : _matrix_c_5_T_15; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 311:30 315:29 320:29]
  wire [63:0] a_tile_v_136_1 = rf_a_tile_v_1_MPORT_136_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] a_tile_v_136_0 = rf_a_tile_v_0_MPORT_136_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_a_5_T_10 = {a_tile_v_136_1,a_tile_v_136_0,128'h0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 325:33]
  wire [63:0] matrix_b_5_tile_v_16_3 = rf_matrix_b_5_tile_v_3_MPORT_16_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_5_tile_v_16_2 = rf_matrix_b_5_tile_v_2_MPORT_16_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_5_tile_v_16_1 = rf_matrix_b_5_tile_v_1_MPORT_16_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_5_tile_v_16_0 = rf_matrix_b_5_tile_v_0_MPORT_16_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_b_5_T_16 = {matrix_b_5_tile_v_16_3,matrix_b_5_tile_v_16_2,matrix_b_5_tile_v_16_1,
    matrix_b_5_tile_v_16_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] matrix_c_5_tile_v_16_3 = rf_matrix_c_5_tile_v_3_MPORT_16_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_5_tile_v_16_2 = rf_matrix_c_5_tile_v_2_MPORT_16_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_5_tile_v_16_1 = rf_matrix_c_5_tile_v_1_MPORT_16_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_5_tile_v_16_0 = rf_matrix_c_5_tile_v_0_MPORT_16_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_c_5_T_16 = {matrix_c_5_tile_v_16_3,matrix_c_5_tile_v_16_2,matrix_c_5_tile_v_16_1,
    matrix_c_5_tile_v_16_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] a_tile_v_137_1 = rf_a_tile_v_1_MPORT_137_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] a_tile_v_137_0 = rf_a_tile_v_0_MPORT_137_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_a_5_T_11 = {a_tile_v_137_1,a_tile_v_137_0,128'h0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 331:33]
  wire [63:0] matrix_b_5_tile_v_17_3 = rf_matrix_b_5_tile_v_3_MPORT_17_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_5_tile_v_17_2 = rf_matrix_b_5_tile_v_2_MPORT_17_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_5_tile_v_17_1 = rf_matrix_b_5_tile_v_1_MPORT_17_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_5_tile_v_17_0 = rf_matrix_b_5_tile_v_0_MPORT_17_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_b_5_T_17 = {matrix_b_5_tile_v_17_3,matrix_b_5_tile_v_17_2,matrix_b_5_tile_v_17_1,
    matrix_b_5_tile_v_17_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] matrix_c_5_tile_v_17_3 = rf_matrix_c_5_tile_v_3_MPORT_17_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_5_tile_v_17_2 = rf_matrix_c_5_tile_v_2_MPORT_17_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_5_tile_v_17_1 = rf_matrix_c_5_tile_v_1_MPORT_17_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_5_tile_v_17_0 = rf_matrix_c_5_tile_v_0_MPORT_17_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_c_5_T_17 = {matrix_c_5_tile_v_17_3,matrix_c_5_tile_v_17_2,matrix_c_5_tile_v_17_1,
    matrix_c_5_tile_v_17_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [255:0] _GEN_8151 = _T_4 ? _matrix_a_5_T_11 : matrix_a_5; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 159:21 296:24 331:27]
  wire [255:0] _GEN_8156 = _T_4 ? _matrix_b_5_T_17 : matrix_b_5; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 160:21 296:24 332:27]
  wire [255:0] _GEN_8161 = _T_4 ? _matrix_c_5_T_17 : matrix_c_5; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 161:21 296:24 333:27]
  wire [255:0] _GEN_8166 = _T_3 ? _matrix_a_5_T_10 : _GEN_8151; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 296:24 325:27]
  wire [255:0] _GEN_8171 = _T_3 ? _matrix_b_5_T_16 : _GEN_8156; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 296:24 326:27]
  wire [255:0] _GEN_8176 = _T_3 ? _matrix_c_5_T_16 : _GEN_8161; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 296:24 327:27]
  wire [255:0] _GEN_8193 = _T_2 ? _GEN_8144 : _GEN_8166; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 296:24]
  wire [255:0] _GEN_8198 = _T_2 ? _GEN_8145 : _GEN_8171; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 296:24]
  wire [255:0] _GEN_8203 = _T_2 ? _GEN_8146 : _GEN_8176; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 296:24]
  wire [255:0] _GEN_8246 = _T_1 ? _GEN_8135 : _GEN_8193; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 296:24]
  wire [255:0] _GEN_8251 = _T_1 ? _GEN_8136 : _GEN_8198; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 296:24]
  wire [255:0] _GEN_8256 = _T_1 ? _GEN_8137 : _GEN_8203; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 296:24]
  wire [63:0] a_tile_v_138_1 = rf_a_tile_v_1_MPORT_138_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] a_tile_v_138_0 = rf_a_tile_v_0_MPORT_138_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_a_5_T_12 = {a_tile_v_138_1,a_tile_v_138_0,128'h0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 342:35]
  wire [63:0] matrix_b_5_tile_v_18_3 = rf_matrix_b_5_tile_v_3_MPORT_18_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_5_tile_v_18_2 = rf_matrix_b_5_tile_v_2_MPORT_18_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_5_tile_v_18_1 = rf_matrix_b_5_tile_v_1_MPORT_18_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_5_tile_v_18_0 = rf_matrix_b_5_tile_v_0_MPORT_18_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_b_5_T_18 = {matrix_b_5_tile_v_18_3,matrix_b_5_tile_v_18_2,matrix_b_5_tile_v_18_1,
    matrix_b_5_tile_v_18_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] matrix_c_5_tile_v_18_3 = rf_matrix_c_5_tile_v_3_MPORT_18_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_5_tile_v_18_2 = rf_matrix_c_5_tile_v_2_MPORT_18_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_5_tile_v_18_1 = rf_matrix_c_5_tile_v_1_MPORT_18_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_5_tile_v_18_0 = rf_matrix_c_5_tile_v_0_MPORT_18_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_c_5_T_18 = {matrix_c_5_tile_v_18_3,matrix_c_5_tile_v_18_2,matrix_c_5_tile_v_18_1,
    matrix_c_5_tile_v_18_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] a_tile_v_139_3 = rf_a_tile_v_3_MPORT_46_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] a_tile_v_139_2 = rf_a_tile_v_2_MPORT_46_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] a_tile_v_139_1 = rf_a_tile_v_1_MPORT_139_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] a_tile_v_139_0 = rf_a_tile_v_0_MPORT_139_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] a_139 = {a_tile_v_139_3,a_tile_v_139_2,a_tile_v_139_1,a_tile_v_139_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] matrix_b_5_tile_v_19_3 = rf_matrix_b_5_tile_v_3_MPORT_19_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_5_tile_v_19_2 = rf_matrix_b_5_tile_v_2_MPORT_19_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_5_tile_v_19_1 = rf_matrix_b_5_tile_v_1_MPORT_19_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_5_tile_v_19_0 = rf_matrix_b_5_tile_v_0_MPORT_19_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_b_5_T_19 = {matrix_b_5_tile_v_19_3,matrix_b_5_tile_v_19_2,matrix_b_5_tile_v_19_1,
    matrix_b_5_tile_v_19_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] matrix_c_5_tile_v_19_3 = rf_matrix_c_5_tile_v_3_MPORT_19_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_5_tile_v_19_2 = rf_matrix_c_5_tile_v_2_MPORT_19_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_5_tile_v_19_1 = rf_matrix_c_5_tile_v_1_MPORT_19_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_5_tile_v_19_0 = rf_matrix_c_5_tile_v_0_MPORT_19_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_c_5_T_19 = {matrix_c_5_tile_v_19_3,matrix_c_5_tile_v_19_2,matrix_c_5_tile_v_19_1,
    matrix_c_5_tile_v_19_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [255:0] _GEN_8323 = io_mixPc ? _matrix_a_5_T_12 : a_139; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 340:30 342:29 347:29]
  wire [255:0] _GEN_8324 = io_mixPc ? _matrix_b_5_T_18 : _matrix_b_5_T_19; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 340:30 343:29 348:29]
  wire [255:0] _GEN_8325 = io_mixPc ? _matrix_c_5_T_18 : _matrix_c_5_T_19; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 340:30 344:29 349:29]
  wire [63:0] a_tile_v_140_1 = rf_a_tile_v_1_MPORT_140_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] a_tile_v_140_0 = rf_a_tile_v_0_MPORT_140_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_a_5_T_13 = {a_tile_v_140_1,a_tile_v_140_0,128'h0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 355:35]
  wire [63:0] matrix_b_5_tile_v_20_3 = rf_matrix_b_5_tile_v_3_MPORT_20_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_5_tile_v_20_2 = rf_matrix_b_5_tile_v_2_MPORT_20_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_5_tile_v_20_1 = rf_matrix_b_5_tile_v_1_MPORT_20_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_5_tile_v_20_0 = rf_matrix_b_5_tile_v_0_MPORT_20_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_b_5_T_20 = {matrix_b_5_tile_v_20_3,matrix_b_5_tile_v_20_2,matrix_b_5_tile_v_20_1,
    matrix_b_5_tile_v_20_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] matrix_c_5_tile_v_20_3 = rf_matrix_c_5_tile_v_3_MPORT_20_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_5_tile_v_20_2 = rf_matrix_c_5_tile_v_2_MPORT_20_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_5_tile_v_20_1 = rf_matrix_c_5_tile_v_1_MPORT_20_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_5_tile_v_20_0 = rf_matrix_c_5_tile_v_0_MPORT_20_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_c_5_T_20 = {matrix_c_5_tile_v_20_3,matrix_c_5_tile_v_20_2,matrix_c_5_tile_v_20_1,
    matrix_c_5_tile_v_20_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] a_tile_v_141_3 = rf_a_tile_v_3_MPORT_47_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] a_tile_v_141_2 = rf_a_tile_v_2_MPORT_47_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] a_tile_v_141_1 = rf_a_tile_v_1_MPORT_141_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] a_tile_v_141_0 = rf_a_tile_v_0_MPORT_141_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] a_141 = {a_tile_v_141_3,a_tile_v_141_2,a_tile_v_141_1,a_tile_v_141_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] matrix_b_5_tile_v_21_3 = rf_matrix_b_5_tile_v_3_MPORT_21_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_5_tile_v_21_2 = rf_matrix_b_5_tile_v_2_MPORT_21_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_5_tile_v_21_1 = rf_matrix_b_5_tile_v_1_MPORT_21_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_5_tile_v_21_0 = rf_matrix_b_5_tile_v_0_MPORT_21_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_b_5_T_21 = {matrix_b_5_tile_v_21_3,matrix_b_5_tile_v_21_2,matrix_b_5_tile_v_21_1,
    matrix_b_5_tile_v_21_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] matrix_c_5_tile_v_21_3 = rf_matrix_c_5_tile_v_3_MPORT_21_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_5_tile_v_21_2 = rf_matrix_c_5_tile_v_2_MPORT_21_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_5_tile_v_21_1 = rf_matrix_c_5_tile_v_1_MPORT_21_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_5_tile_v_21_0 = rf_matrix_c_5_tile_v_0_MPORT_21_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_c_5_T_21 = {matrix_c_5_tile_v_21_3,matrix_c_5_tile_v_21_2,matrix_c_5_tile_v_21_1,
    matrix_c_5_tile_v_21_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [255:0] _GEN_8332 = io_mixPc ? _matrix_a_5_T_13 : a_141; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 353:30 355:29 360:29]
  wire [255:0] _GEN_8333 = io_mixPc ? _matrix_b_5_T_20 : _matrix_b_5_T_21; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 353:30 356:29 361:29]
  wire [255:0] _GEN_8334 = io_mixPc ? _matrix_c_5_T_20 : _matrix_c_5_T_21; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 353:30 357:29 362:29]
  wire [63:0] a_tile_v_142_1 = rf_a_tile_v_1_MPORT_142_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] a_tile_v_142_0 = rf_a_tile_v_0_MPORT_142_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_a_5_T_14 = {a_tile_v_142_1,a_tile_v_142_0,128'h0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 367:33]
  wire [63:0] matrix_b_5_tile_v_22_3 = rf_matrix_b_5_tile_v_3_MPORT_22_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_5_tile_v_22_2 = rf_matrix_b_5_tile_v_2_MPORT_22_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_5_tile_v_22_1 = rf_matrix_b_5_tile_v_1_MPORT_22_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_5_tile_v_22_0 = rf_matrix_b_5_tile_v_0_MPORT_22_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_b_5_T_22 = {matrix_b_5_tile_v_22_3,matrix_b_5_tile_v_22_2,matrix_b_5_tile_v_22_1,
    matrix_b_5_tile_v_22_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] matrix_c_5_tile_v_22_3 = rf_matrix_c_5_tile_v_3_MPORT_22_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_5_tile_v_22_2 = rf_matrix_c_5_tile_v_2_MPORT_22_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_5_tile_v_22_1 = rf_matrix_c_5_tile_v_1_MPORT_22_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_5_tile_v_22_0 = rf_matrix_c_5_tile_v_0_MPORT_22_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_c_5_T_22 = {matrix_c_5_tile_v_22_3,matrix_c_5_tile_v_22_2,matrix_c_5_tile_v_22_1,
    matrix_c_5_tile_v_22_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] a_tile_v_143_1 = rf_a_tile_v_1_MPORT_143_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] a_tile_v_143_0 = rf_a_tile_v_0_MPORT_143_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_a_5_T_15 = {a_tile_v_143_1,a_tile_v_143_0,128'h0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 373:33]
  wire [63:0] matrix_b_5_tile_v_23_3 = rf_matrix_b_5_tile_v_3_MPORT_23_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_5_tile_v_23_2 = rf_matrix_b_5_tile_v_2_MPORT_23_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_5_tile_v_23_1 = rf_matrix_b_5_tile_v_1_MPORT_23_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_5_tile_v_23_0 = rf_matrix_b_5_tile_v_0_MPORT_23_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_b_5_T_23 = {matrix_b_5_tile_v_23_3,matrix_b_5_tile_v_23_2,matrix_b_5_tile_v_23_1,
    matrix_b_5_tile_v_23_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] matrix_c_5_tile_v_23_3 = rf_matrix_c_5_tile_v_3_MPORT_23_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_5_tile_v_23_2 = rf_matrix_c_5_tile_v_2_MPORT_23_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_5_tile_v_23_1 = rf_matrix_c_5_tile_v_1_MPORT_23_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_5_tile_v_23_0 = rf_matrix_c_5_tile_v_0_MPORT_23_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_c_5_T_23 = {matrix_c_5_tile_v_23_3,matrix_c_5_tile_v_23_2,matrix_c_5_tile_v_23_1,
    matrix_c_5_tile_v_23_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [255:0] _GEN_8339 = _T_4 ? _matrix_a_5_T_15 : matrix_a_5; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 159:21 338:24 373:27]
  wire [255:0] _GEN_8344 = _T_4 ? _matrix_b_5_T_23 : matrix_b_5; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 160:21 338:24 374:27]
  wire [255:0] _GEN_8349 = _T_4 ? _matrix_c_5_T_23 : matrix_c_5; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 161:21 338:24 375:27]
  wire [255:0] _GEN_8354 = _T_3 ? _matrix_a_5_T_14 : _GEN_8339; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 338:24 367:27]
  wire [255:0] _GEN_8359 = _T_3 ? _matrix_b_5_T_22 : _GEN_8344; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 338:24 368:27]
  wire [255:0] _GEN_8364 = _T_3 ? _matrix_c_5_T_22 : _GEN_8349; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 338:24 369:27]
  wire [255:0] _GEN_8381 = _T_2 ? _GEN_8332 : _GEN_8354; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 338:24]
  wire [255:0] _GEN_8386 = _T_2 ? _GEN_8333 : _GEN_8359; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 338:24]
  wire [255:0] _GEN_8391 = _T_2 ? _GEN_8334 : _GEN_8364; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 338:24]
  wire [255:0] _GEN_8434 = _T_1 ? _GEN_8323 : _GEN_8381; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 338:24]
  wire [255:0] _GEN_8439 = _T_1 ? _GEN_8324 : _GEN_8386; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 338:24]
  wire [255:0] _GEN_8444 = _T_1 ? _GEN_8325 : _GEN_8391; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 338:24]
  wire [255:0] _GEN_8513 = 2'h3 == set ? _GEN_8434 : matrix_a_5; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 210:18 159:21]
  wire [255:0] _GEN_8518 = 2'h3 == set ? _GEN_8439 : matrix_b_5; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 210:18 160:21]
  wire [255:0] _GEN_8523 = 2'h3 == set ? _GEN_8444 : matrix_c_5; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 210:18 161:21]
  wire [63:0] a_tile_v_144_1 = rf_a_tile_v_1_MPORT_144_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] a_tile_v_144_0 = rf_a_tile_v_0_MPORT_144_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_a_6_T = {a_tile_v_144_1,a_tile_v_144_0,128'h0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 216:35]
  wire [63:0] matrix_b_6_tile_v__3 = rf_matrix_b_6_tile_v_3_MPORT_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_6_tile_v__2 = rf_matrix_b_6_tile_v_2_MPORT_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_6_tile_v__1 = rf_matrix_b_6_tile_v_1_MPORT_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_6_tile_v__0 = rf_matrix_b_6_tile_v_0_MPORT_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_b_6_T = {matrix_b_6_tile_v__3,matrix_b_6_tile_v__2,matrix_b_6_tile_v__1,matrix_b_6_tile_v__0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] matrix_c_6_tile_v__3 = rf_matrix_c_6_tile_v_3_MPORT_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_6_tile_v__2 = rf_matrix_c_6_tile_v_2_MPORT_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_6_tile_v__1 = rf_matrix_c_6_tile_v_1_MPORT_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_6_tile_v__0 = rf_matrix_c_6_tile_v_0_MPORT_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_c_6_T = {matrix_c_6_tile_v__3,matrix_c_6_tile_v__2,matrix_c_6_tile_v__1,matrix_c_6_tile_v__0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] a_tile_v_145_3 = rf_a_tile_v_3_MPORT_48_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] a_tile_v_145_2 = rf_a_tile_v_2_MPORT_48_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] a_tile_v_145_1 = rf_a_tile_v_1_MPORT_145_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] a_tile_v_145_0 = rf_a_tile_v_0_MPORT_145_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] a_145 = {a_tile_v_145_3,a_tile_v_145_2,a_tile_v_145_1,a_tile_v_145_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] matrix_b_6_tile_v_1_3 = rf_matrix_b_6_tile_v_3_MPORT_1_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_6_tile_v_1_2 = rf_matrix_b_6_tile_v_2_MPORT_1_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_6_tile_v_1_1 = rf_matrix_b_6_tile_v_1_MPORT_1_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_6_tile_v_1_0 = rf_matrix_b_6_tile_v_0_MPORT_1_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_b_6_T_1 = {matrix_b_6_tile_v_1_3,matrix_b_6_tile_v_1_2,matrix_b_6_tile_v_1_1,
    matrix_b_6_tile_v_1_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] matrix_c_6_tile_v_1_3 = rf_matrix_c_6_tile_v_3_MPORT_1_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_6_tile_v_1_2 = rf_matrix_c_6_tile_v_2_MPORT_1_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_6_tile_v_1_1 = rf_matrix_c_6_tile_v_1_MPORT_1_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_6_tile_v_1_0 = rf_matrix_c_6_tile_v_0_MPORT_1_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_c_6_T_1 = {matrix_c_6_tile_v_1_3,matrix_c_6_tile_v_1_2,matrix_c_6_tile_v_1_1,
    matrix_c_6_tile_v_1_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] a_tile_v_146_1 = rf_a_tile_v_1_MPORT_146_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] a_tile_v_146_0 = rf_a_tile_v_0_MPORT_146_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_a_6_T_1 = {a_tile_v_146_1,a_tile_v_146_0,128'h0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 229:35]
  wire [63:0] matrix_b_6_tile_v_2_3 = rf_matrix_b_6_tile_v_3_MPORT_2_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_6_tile_v_2_2 = rf_matrix_b_6_tile_v_2_MPORT_2_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_6_tile_v_2_1 = rf_matrix_b_6_tile_v_1_MPORT_2_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_6_tile_v_2_0 = rf_matrix_b_6_tile_v_0_MPORT_2_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_b_6_T_2 = {matrix_b_6_tile_v_2_3,matrix_b_6_tile_v_2_2,matrix_b_6_tile_v_2_1,
    matrix_b_6_tile_v_2_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] matrix_c_6_tile_v_2_3 = rf_matrix_c_6_tile_v_3_MPORT_2_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_6_tile_v_2_2 = rf_matrix_c_6_tile_v_2_MPORT_2_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_6_tile_v_2_1 = rf_matrix_c_6_tile_v_1_MPORT_2_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_6_tile_v_2_0 = rf_matrix_c_6_tile_v_0_MPORT_2_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_c_6_T_2 = {matrix_c_6_tile_v_2_3,matrix_c_6_tile_v_2_2,matrix_c_6_tile_v_2_1,
    matrix_c_6_tile_v_2_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] a_tile_v_147_3 = rf_a_tile_v_3_MPORT_49_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] a_tile_v_147_2 = rf_a_tile_v_2_MPORT_49_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] a_tile_v_147_1 = rf_a_tile_v_1_MPORT_147_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] a_tile_v_147_0 = rf_a_tile_v_0_MPORT_147_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] a_147 = {a_tile_v_147_3,a_tile_v_147_2,a_tile_v_147_1,a_tile_v_147_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] matrix_b_6_tile_v_3_3 = rf_matrix_b_6_tile_v_3_MPORT_3_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_6_tile_v_3_2 = rf_matrix_b_6_tile_v_2_MPORT_3_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_6_tile_v_3_1 = rf_matrix_b_6_tile_v_1_MPORT_3_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_6_tile_v_3_0 = rf_matrix_b_6_tile_v_0_MPORT_3_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_b_6_T_3 = {matrix_b_6_tile_v_3_3,matrix_b_6_tile_v_3_2,matrix_b_6_tile_v_3_1,
    matrix_b_6_tile_v_3_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] matrix_c_6_tile_v_3_3 = rf_matrix_c_6_tile_v_3_MPORT_3_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_6_tile_v_3_2 = rf_matrix_c_6_tile_v_2_MPORT_3_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_6_tile_v_3_1 = rf_matrix_c_6_tile_v_1_MPORT_3_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_6_tile_v_3_0 = rf_matrix_c_6_tile_v_0_MPORT_3_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_c_6_T_3 = {matrix_c_6_tile_v_3_3,matrix_c_6_tile_v_3_2,matrix_c_6_tile_v_3_1,
    matrix_c_6_tile_v_3_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [255:0] _GEN_9300 = io_mixPc ? _matrix_a_6_T_1 : a_147; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 227:30 229:29 234:29]
  wire [255:0] _GEN_9301 = io_mixPc ? _matrix_b_6_T_2 : _matrix_b_6_T_3; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 227:30 230:29 235:29]
  wire [255:0] _GEN_9306 = io_mixPc ? _matrix_c_6_T_2 : _matrix_c_6_T_3; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 227:30 231:29 236:29]
  wire [63:0] a_tile_v_148_1 = rf_a_tile_v_1_MPORT_148_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] a_tile_v_148_0 = rf_a_tile_v_0_MPORT_148_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_a_6_T_2 = {a_tile_v_148_1,a_tile_v_148_0,128'h0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 241:33]
  wire [63:0] matrix_b_6_tile_v_4_3 = rf_matrix_b_6_tile_v_3_MPORT_4_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_6_tile_v_4_2 = rf_matrix_b_6_tile_v_2_MPORT_4_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_6_tile_v_4_1 = rf_matrix_b_6_tile_v_1_MPORT_4_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_6_tile_v_4_0 = rf_matrix_b_6_tile_v_0_MPORT_4_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_b_6_T_4 = {matrix_b_6_tile_v_4_3,matrix_b_6_tile_v_4_2,matrix_b_6_tile_v_4_1,
    matrix_b_6_tile_v_4_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] matrix_c_6_tile_v_4_3 = rf_matrix_c_6_tile_v_3_MPORT_4_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_6_tile_v_4_2 = rf_matrix_c_6_tile_v_2_MPORT_4_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_6_tile_v_4_1 = rf_matrix_c_6_tile_v_1_MPORT_4_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_6_tile_v_4_0 = rf_matrix_c_6_tile_v_0_MPORT_4_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_c_6_T_4 = {matrix_c_6_tile_v_4_3,matrix_c_6_tile_v_4_2,matrix_c_6_tile_v_4_1,
    matrix_c_6_tile_v_4_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] a_tile_v_149_1 = rf_a_tile_v_1_MPORT_149_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] a_tile_v_149_0 = rf_a_tile_v_0_MPORT_149_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_a_6_T_3 = {a_tile_v_149_1,a_tile_v_149_0,128'h0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 247:33]
  wire [63:0] matrix_b_6_tile_v_5_3 = rf_matrix_b_6_tile_v_3_MPORT_5_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_6_tile_v_5_2 = rf_matrix_b_6_tile_v_2_MPORT_5_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_6_tile_v_5_1 = rf_matrix_b_6_tile_v_1_MPORT_5_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_6_tile_v_5_0 = rf_matrix_b_6_tile_v_0_MPORT_5_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_b_6_T_5 = {matrix_b_6_tile_v_5_3,matrix_b_6_tile_v_5_2,matrix_b_6_tile_v_5_1,
    matrix_b_6_tile_v_5_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] matrix_c_6_tile_v_5_3 = rf_matrix_c_6_tile_v_3_MPORT_5_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_6_tile_v_5_2 = rf_matrix_c_6_tile_v_2_MPORT_5_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_6_tile_v_5_1 = rf_matrix_c_6_tile_v_1_MPORT_5_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_6_tile_v_5_0 = rf_matrix_c_6_tile_v_0_MPORT_5_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_c_6_T_5 = {matrix_c_6_tile_v_5_3,matrix_c_6_tile_v_5_2,matrix_c_6_tile_v_5_1,
    matrix_c_6_tile_v_5_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [255:0] _GEN_9315 = 2'h3 == step ? _matrix_a_6_T_3 : matrix_a_6; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 159:21 212:23 247:27]
  wire [255:0] _GEN_9320 = 2'h3 == step ? _matrix_b_6_T_5 : matrix_b_6; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 160:21 212:23 248:27]
  wire [255:0] _GEN_9325 = 2'h3 == step ? _matrix_c_6_T_5 : matrix_c_6; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 161:21 212:23 249:27]
  wire [255:0] _GEN_9330 = 2'h2 == step ? _matrix_a_6_T_2 : _GEN_9315; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 212:23 241:27]
  wire [255:0] _GEN_9335 = 2'h2 == step ? _matrix_b_6_T_4 : _GEN_9320; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 212:23 242:27]
  wire [255:0] _GEN_9340 = 2'h2 == step ? _matrix_c_6_T_4 : _GEN_9325; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 212:23 243:27]
  wire [63:0] a_tile_v_150_1 = rf_a_tile_v_1_MPORT_150_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] a_tile_v_150_0 = rf_a_tile_v_0_MPORT_150_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_a_6_T_4 = {a_tile_v_150_1,a_tile_v_150_0,128'h0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 258:35]
  wire [63:0] matrix_b_6_tile_v_6_3 = rf_matrix_b_6_tile_v_3_MPORT_6_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_6_tile_v_6_2 = rf_matrix_b_6_tile_v_2_MPORT_6_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_6_tile_v_6_1 = rf_matrix_b_6_tile_v_1_MPORT_6_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_6_tile_v_6_0 = rf_matrix_b_6_tile_v_0_MPORT_6_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_b_6_T_6 = {matrix_b_6_tile_v_6_3,matrix_b_6_tile_v_6_2,matrix_b_6_tile_v_6_1,
    matrix_b_6_tile_v_6_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] matrix_c_6_tile_v_6_3 = rf_matrix_c_6_tile_v_3_MPORT_6_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_6_tile_v_6_2 = rf_matrix_c_6_tile_v_2_MPORT_6_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_6_tile_v_6_1 = rf_matrix_c_6_tile_v_1_MPORT_6_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_6_tile_v_6_0 = rf_matrix_c_6_tile_v_0_MPORT_6_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_c_6_T_6 = {matrix_c_6_tile_v_6_3,matrix_c_6_tile_v_6_2,matrix_c_6_tile_v_6_1,
    matrix_c_6_tile_v_6_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] a_tile_v_151_3 = rf_a_tile_v_3_MPORT_50_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] a_tile_v_151_2 = rf_a_tile_v_2_MPORT_50_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] a_tile_v_151_1 = rf_a_tile_v_1_MPORT_151_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] a_tile_v_151_0 = rf_a_tile_v_0_MPORT_151_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] a_151 = {a_tile_v_151_3,a_tile_v_151_2,a_tile_v_151_1,a_tile_v_151_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] matrix_b_6_tile_v_7_3 = rf_matrix_b_6_tile_v_3_MPORT_7_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_6_tile_v_7_2 = rf_matrix_b_6_tile_v_2_MPORT_7_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_6_tile_v_7_1 = rf_matrix_b_6_tile_v_1_MPORT_7_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_6_tile_v_7_0 = rf_matrix_b_6_tile_v_0_MPORT_7_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_b_6_T_7 = {matrix_b_6_tile_v_7_3,matrix_b_6_tile_v_7_2,matrix_b_6_tile_v_7_1,
    matrix_b_6_tile_v_7_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] matrix_c_6_tile_v_7_3 = rf_matrix_c_6_tile_v_3_MPORT_7_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_6_tile_v_7_2 = rf_matrix_c_6_tile_v_2_MPORT_7_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_6_tile_v_7_1 = rf_matrix_c_6_tile_v_1_MPORT_7_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_6_tile_v_7_0 = rf_matrix_c_6_tile_v_0_MPORT_7_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_c_6_T_7 = {matrix_c_6_tile_v_7_3,matrix_c_6_tile_v_7_2,matrix_c_6_tile_v_7_1,
    matrix_c_6_tile_v_7_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [255:0] _GEN_9485 = io_mixPc ? _matrix_a_6_T_4 : a_151; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 256:30 258:29 263:29]
  wire [255:0] _GEN_9490 = io_mixPc ? _matrix_b_6_T_6 : _matrix_b_6_T_7; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 256:30 259:29 264:29]
  wire [255:0] _GEN_9491 = io_mixPc ? _matrix_c_6_T_6 : _matrix_c_6_T_7; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 256:30 260:29 265:29]
  wire [63:0] a_tile_v_152_1 = rf_a_tile_v_1_MPORT_152_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] a_tile_v_152_0 = rf_a_tile_v_0_MPORT_152_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_a_6_T_5 = {a_tile_v_152_1,a_tile_v_152_0,128'h0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 271:35]
  wire [63:0] matrix_b_6_tile_v_8_3 = rf_matrix_b_6_tile_v_3_MPORT_8_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_6_tile_v_8_2 = rf_matrix_b_6_tile_v_2_MPORT_8_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_6_tile_v_8_1 = rf_matrix_b_6_tile_v_1_MPORT_8_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_6_tile_v_8_0 = rf_matrix_b_6_tile_v_0_MPORT_8_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_b_6_T_8 = {matrix_b_6_tile_v_8_3,matrix_b_6_tile_v_8_2,matrix_b_6_tile_v_8_1,
    matrix_b_6_tile_v_8_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] matrix_c_6_tile_v_8_3 = rf_matrix_c_6_tile_v_3_MPORT_8_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_6_tile_v_8_2 = rf_matrix_c_6_tile_v_2_MPORT_8_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_6_tile_v_8_1 = rf_matrix_c_6_tile_v_1_MPORT_8_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_6_tile_v_8_0 = rf_matrix_c_6_tile_v_0_MPORT_8_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_c_6_T_8 = {matrix_c_6_tile_v_8_3,matrix_c_6_tile_v_8_2,matrix_c_6_tile_v_8_1,
    matrix_c_6_tile_v_8_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] a_tile_v_153_3 = rf_a_tile_v_3_MPORT_51_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] a_tile_v_153_2 = rf_a_tile_v_2_MPORT_51_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] a_tile_v_153_1 = rf_a_tile_v_1_MPORT_153_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] a_tile_v_153_0 = rf_a_tile_v_0_MPORT_153_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] a_153 = {a_tile_v_153_3,a_tile_v_153_2,a_tile_v_153_1,a_tile_v_153_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] matrix_b_6_tile_v_9_3 = rf_matrix_b_6_tile_v_3_MPORT_9_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_6_tile_v_9_2 = rf_matrix_b_6_tile_v_2_MPORT_9_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_6_tile_v_9_1 = rf_matrix_b_6_tile_v_1_MPORT_9_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_6_tile_v_9_0 = rf_matrix_b_6_tile_v_0_MPORT_9_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_b_6_T_9 = {matrix_b_6_tile_v_9_3,matrix_b_6_tile_v_9_2,matrix_b_6_tile_v_9_1,
    matrix_b_6_tile_v_9_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] matrix_c_6_tile_v_9_3 = rf_matrix_c_6_tile_v_3_MPORT_9_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_6_tile_v_9_2 = rf_matrix_c_6_tile_v_2_MPORT_9_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_6_tile_v_9_1 = rf_matrix_c_6_tile_v_1_MPORT_9_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_6_tile_v_9_0 = rf_matrix_c_6_tile_v_0_MPORT_9_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_c_6_T_9 = {matrix_c_6_tile_v_9_3,matrix_c_6_tile_v_9_2,matrix_c_6_tile_v_9_1,
    matrix_c_6_tile_v_9_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [255:0] _GEN_9496 = io_mixPc ? _matrix_a_6_T_5 : a_153; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 269:30 271:29 276:29]
  wire [255:0] _GEN_9497 = io_mixPc ? _matrix_b_6_T_8 : _matrix_b_6_T_9; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 269:30 272:29 277:29]
  wire [255:0] _GEN_9498 = io_mixPc ? _matrix_c_6_T_8 : _matrix_c_6_T_9; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 269:30 273:29 278:29]
  wire [63:0] a_tile_v_154_1 = rf_a_tile_v_1_MPORT_154_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] a_tile_v_154_0 = rf_a_tile_v_0_MPORT_154_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_a_6_T_6 = {a_tile_v_154_1,a_tile_v_154_0,128'h0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 283:33]
  wire [63:0] matrix_b_6_tile_v_10_3 = rf_matrix_b_6_tile_v_3_MPORT_10_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_6_tile_v_10_2 = rf_matrix_b_6_tile_v_2_MPORT_10_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_6_tile_v_10_1 = rf_matrix_b_6_tile_v_1_MPORT_10_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_6_tile_v_10_0 = rf_matrix_b_6_tile_v_0_MPORT_10_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_b_6_T_10 = {matrix_b_6_tile_v_10_3,matrix_b_6_tile_v_10_2,matrix_b_6_tile_v_10_1,
    matrix_b_6_tile_v_10_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] matrix_c_6_tile_v_10_3 = rf_matrix_c_6_tile_v_3_MPORT_10_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_6_tile_v_10_2 = rf_matrix_c_6_tile_v_2_MPORT_10_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_6_tile_v_10_1 = rf_matrix_c_6_tile_v_1_MPORT_10_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_6_tile_v_10_0 = rf_matrix_c_6_tile_v_0_MPORT_10_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_c_6_T_10 = {matrix_c_6_tile_v_10_3,matrix_c_6_tile_v_10_2,matrix_c_6_tile_v_10_1,
    matrix_c_6_tile_v_10_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] a_tile_v_155_1 = rf_a_tile_v_1_MPORT_155_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] a_tile_v_155_0 = rf_a_tile_v_0_MPORT_155_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_a_6_T_7 = {a_tile_v_155_1,a_tile_v_155_0,128'h0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 289:33]
  wire [63:0] matrix_b_6_tile_v_11_3 = rf_matrix_b_6_tile_v_3_MPORT_11_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_6_tile_v_11_2 = rf_matrix_b_6_tile_v_2_MPORT_11_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_6_tile_v_11_1 = rf_matrix_b_6_tile_v_1_MPORT_11_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_6_tile_v_11_0 = rf_matrix_b_6_tile_v_0_MPORT_11_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_b_6_T_11 = {matrix_b_6_tile_v_11_3,matrix_b_6_tile_v_11_2,matrix_b_6_tile_v_11_1,
    matrix_b_6_tile_v_11_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] matrix_c_6_tile_v_11_3 = rf_matrix_c_6_tile_v_3_MPORT_11_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_6_tile_v_11_2 = rf_matrix_c_6_tile_v_2_MPORT_11_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_6_tile_v_11_1 = rf_matrix_c_6_tile_v_1_MPORT_11_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_6_tile_v_11_0 = rf_matrix_c_6_tile_v_0_MPORT_11_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_c_6_T_11 = {matrix_c_6_tile_v_11_3,matrix_c_6_tile_v_11_2,matrix_c_6_tile_v_11_1,
    matrix_c_6_tile_v_11_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [255:0] _GEN_9503 = _T_4 ? _matrix_a_6_T_7 : matrix_a_6; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 159:21 254:24 289:27]
  wire [255:0] _GEN_9508 = _T_4 ? _matrix_b_6_T_11 : matrix_b_6; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 160:21 254:24 290:27]
  wire [255:0] _GEN_9513 = _T_4 ? _matrix_c_6_T_11 : matrix_c_6; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 161:21 254:24 291:27]
  wire [255:0] _GEN_9518 = _T_3 ? _matrix_a_6_T_6 : _GEN_9503; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 254:24 283:27]
  wire [255:0] _GEN_9523 = _T_3 ? _matrix_b_6_T_10 : _GEN_9508; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 254:24 284:27]
  wire [255:0] _GEN_9528 = _T_3 ? _matrix_c_6_T_10 : _GEN_9513; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 254:24 285:27]
  wire [255:0] _GEN_9545 = _T_2 ? _GEN_9496 : _GEN_9518; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 254:24]
  wire [255:0] _GEN_9550 = _T_2 ? _GEN_9497 : _GEN_9523; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 254:24]
  wire [255:0] _GEN_9555 = _T_2 ? _GEN_9498 : _GEN_9528; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 254:24]
  wire [63:0] a_tile_v_156_1 = rf_a_tile_v_1_MPORT_156_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] a_tile_v_156_0 = rf_a_tile_v_0_MPORT_156_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_a_6_T_8 = {a_tile_v_156_1,a_tile_v_156_0,128'h0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 300:35]
  wire [63:0] matrix_b_6_tile_v_12_3 = rf_matrix_b_6_tile_v_3_MPORT_12_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_6_tile_v_12_2 = rf_matrix_b_6_tile_v_2_MPORT_12_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_6_tile_v_12_1 = rf_matrix_b_6_tile_v_1_MPORT_12_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_6_tile_v_12_0 = rf_matrix_b_6_tile_v_0_MPORT_12_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_b_6_T_12 = {matrix_b_6_tile_v_12_3,matrix_b_6_tile_v_12_2,matrix_b_6_tile_v_12_1,
    matrix_b_6_tile_v_12_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] matrix_c_6_tile_v_12_3 = rf_matrix_c_6_tile_v_3_MPORT_12_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_6_tile_v_12_2 = rf_matrix_c_6_tile_v_2_MPORT_12_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_6_tile_v_12_1 = rf_matrix_c_6_tile_v_1_MPORT_12_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_6_tile_v_12_0 = rf_matrix_c_6_tile_v_0_MPORT_12_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_c_6_T_12 = {matrix_c_6_tile_v_12_3,matrix_c_6_tile_v_12_2,matrix_c_6_tile_v_12_1,
    matrix_c_6_tile_v_12_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] a_tile_v_157_3 = rf_a_tile_v_3_MPORT_52_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] a_tile_v_157_2 = rf_a_tile_v_2_MPORT_52_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] a_tile_v_157_1 = rf_a_tile_v_1_MPORT_157_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] a_tile_v_157_0 = rf_a_tile_v_0_MPORT_157_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] a_157 = {a_tile_v_157_3,a_tile_v_157_2,a_tile_v_157_1,a_tile_v_157_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] matrix_b_6_tile_v_13_3 = rf_matrix_b_6_tile_v_3_MPORT_13_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_6_tile_v_13_2 = rf_matrix_b_6_tile_v_2_MPORT_13_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_6_tile_v_13_1 = rf_matrix_b_6_tile_v_1_MPORT_13_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_6_tile_v_13_0 = rf_matrix_b_6_tile_v_0_MPORT_13_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_b_6_T_13 = {matrix_b_6_tile_v_13_3,matrix_b_6_tile_v_13_2,matrix_b_6_tile_v_13_1,
    matrix_b_6_tile_v_13_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] matrix_c_6_tile_v_13_3 = rf_matrix_c_6_tile_v_3_MPORT_13_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_6_tile_v_13_2 = rf_matrix_c_6_tile_v_2_MPORT_13_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_6_tile_v_13_1 = rf_matrix_c_6_tile_v_1_MPORT_13_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_6_tile_v_13_0 = rf_matrix_c_6_tile_v_0_MPORT_13_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_c_6_T_13 = {matrix_c_6_tile_v_13_3,matrix_c_6_tile_v_13_2,matrix_c_6_tile_v_13_1,
    matrix_c_6_tile_v_13_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [255:0] _GEN_9673 = io_mixPc ? _matrix_a_6_T_8 : a_157; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 298:30 300:29 305:29]
  wire [255:0] _GEN_9678 = io_mixPc ? _matrix_b_6_T_12 : _matrix_b_6_T_13; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 298:30 301:29 306:29]
  wire [255:0] _GEN_9679 = io_mixPc ? _matrix_c_6_T_12 : _matrix_c_6_T_13; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 298:30 302:29 307:29]
  wire [63:0] a_tile_v_158_1 = rf_a_tile_v_1_MPORT_158_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] a_tile_v_158_0 = rf_a_tile_v_0_MPORT_158_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_a_6_T_9 = {a_tile_v_158_1,a_tile_v_158_0,128'h0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 313:35]
  wire [63:0] matrix_b_6_tile_v_14_3 = rf_matrix_b_6_tile_v_3_MPORT_14_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_6_tile_v_14_2 = rf_matrix_b_6_tile_v_2_MPORT_14_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_6_tile_v_14_1 = rf_matrix_b_6_tile_v_1_MPORT_14_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_6_tile_v_14_0 = rf_matrix_b_6_tile_v_0_MPORT_14_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_b_6_T_14 = {matrix_b_6_tile_v_14_3,matrix_b_6_tile_v_14_2,matrix_b_6_tile_v_14_1,
    matrix_b_6_tile_v_14_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] matrix_c_6_tile_v_14_3 = rf_matrix_c_6_tile_v_3_MPORT_14_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_6_tile_v_14_2 = rf_matrix_c_6_tile_v_2_MPORT_14_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_6_tile_v_14_1 = rf_matrix_c_6_tile_v_1_MPORT_14_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_6_tile_v_14_0 = rf_matrix_c_6_tile_v_0_MPORT_14_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_c_6_T_14 = {matrix_c_6_tile_v_14_3,matrix_c_6_tile_v_14_2,matrix_c_6_tile_v_14_1,
    matrix_c_6_tile_v_14_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] a_tile_v_159_3 = rf_a_tile_v_3_MPORT_53_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] a_tile_v_159_2 = rf_a_tile_v_2_MPORT_53_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] a_tile_v_159_1 = rf_a_tile_v_1_MPORT_159_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] a_tile_v_159_0 = rf_a_tile_v_0_MPORT_159_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] a_159 = {a_tile_v_159_3,a_tile_v_159_2,a_tile_v_159_1,a_tile_v_159_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] matrix_b_6_tile_v_15_3 = rf_matrix_b_6_tile_v_3_MPORT_15_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_6_tile_v_15_2 = rf_matrix_b_6_tile_v_2_MPORT_15_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_6_tile_v_15_1 = rf_matrix_b_6_tile_v_1_MPORT_15_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_6_tile_v_15_0 = rf_matrix_b_6_tile_v_0_MPORT_15_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_b_6_T_15 = {matrix_b_6_tile_v_15_3,matrix_b_6_tile_v_15_2,matrix_b_6_tile_v_15_1,
    matrix_b_6_tile_v_15_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] matrix_c_6_tile_v_15_3 = rf_matrix_c_6_tile_v_3_MPORT_15_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_6_tile_v_15_2 = rf_matrix_c_6_tile_v_2_MPORT_15_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_6_tile_v_15_1 = rf_matrix_c_6_tile_v_1_MPORT_15_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_6_tile_v_15_0 = rf_matrix_c_6_tile_v_0_MPORT_15_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_c_6_T_15 = {matrix_c_6_tile_v_15_3,matrix_c_6_tile_v_15_2,matrix_c_6_tile_v_15_1,
    matrix_c_6_tile_v_15_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [255:0] _GEN_9684 = io_mixPc ? _matrix_a_6_T_9 : a_159; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 311:30 313:29 318:29]
  wire [255:0] _GEN_9685 = io_mixPc ? _matrix_b_6_T_14 : _matrix_b_6_T_15; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 311:30 314:29 319:29]
  wire [255:0] _GEN_9686 = io_mixPc ? _matrix_c_6_T_14 : _matrix_c_6_T_15; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 311:30 315:29 320:29]
  wire [63:0] a_tile_v_160_1 = rf_a_tile_v_1_MPORT_160_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] a_tile_v_160_0 = rf_a_tile_v_0_MPORT_160_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_a_6_T_10 = {a_tile_v_160_1,a_tile_v_160_0,128'h0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 325:33]
  wire [63:0] matrix_b_6_tile_v_16_3 = rf_matrix_b_6_tile_v_3_MPORT_16_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_6_tile_v_16_2 = rf_matrix_b_6_tile_v_2_MPORT_16_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_6_tile_v_16_1 = rf_matrix_b_6_tile_v_1_MPORT_16_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_6_tile_v_16_0 = rf_matrix_b_6_tile_v_0_MPORT_16_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_b_6_T_16 = {matrix_b_6_tile_v_16_3,matrix_b_6_tile_v_16_2,matrix_b_6_tile_v_16_1,
    matrix_b_6_tile_v_16_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] matrix_c_6_tile_v_16_3 = rf_matrix_c_6_tile_v_3_MPORT_16_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_6_tile_v_16_2 = rf_matrix_c_6_tile_v_2_MPORT_16_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_6_tile_v_16_1 = rf_matrix_c_6_tile_v_1_MPORT_16_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_6_tile_v_16_0 = rf_matrix_c_6_tile_v_0_MPORT_16_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_c_6_T_16 = {matrix_c_6_tile_v_16_3,matrix_c_6_tile_v_16_2,matrix_c_6_tile_v_16_1,
    matrix_c_6_tile_v_16_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] a_tile_v_161_1 = rf_a_tile_v_1_MPORT_161_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] a_tile_v_161_0 = rf_a_tile_v_0_MPORT_161_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_a_6_T_11 = {a_tile_v_161_1,a_tile_v_161_0,128'h0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 331:33]
  wire [63:0] matrix_b_6_tile_v_17_3 = rf_matrix_b_6_tile_v_3_MPORT_17_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_6_tile_v_17_2 = rf_matrix_b_6_tile_v_2_MPORT_17_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_6_tile_v_17_1 = rf_matrix_b_6_tile_v_1_MPORT_17_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_6_tile_v_17_0 = rf_matrix_b_6_tile_v_0_MPORT_17_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_b_6_T_17 = {matrix_b_6_tile_v_17_3,matrix_b_6_tile_v_17_2,matrix_b_6_tile_v_17_1,
    matrix_b_6_tile_v_17_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] matrix_c_6_tile_v_17_3 = rf_matrix_c_6_tile_v_3_MPORT_17_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_6_tile_v_17_2 = rf_matrix_c_6_tile_v_2_MPORT_17_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_6_tile_v_17_1 = rf_matrix_c_6_tile_v_1_MPORT_17_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_6_tile_v_17_0 = rf_matrix_c_6_tile_v_0_MPORT_17_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_c_6_T_17 = {matrix_c_6_tile_v_17_3,matrix_c_6_tile_v_17_2,matrix_c_6_tile_v_17_1,
    matrix_c_6_tile_v_17_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [255:0] _GEN_9691 = _T_4 ? _matrix_a_6_T_11 : matrix_a_6; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 159:21 296:24 331:27]
  wire [255:0] _GEN_9696 = _T_4 ? _matrix_b_6_T_17 : matrix_b_6; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 160:21 296:24 332:27]
  wire [255:0] _GEN_9701 = _T_4 ? _matrix_c_6_T_17 : matrix_c_6; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 161:21 296:24 333:27]
  wire [255:0] _GEN_9706 = _T_3 ? _matrix_a_6_T_10 : _GEN_9691; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 296:24 325:27]
  wire [255:0] _GEN_9711 = _T_3 ? _matrix_b_6_T_16 : _GEN_9696; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 296:24 326:27]
  wire [255:0] _GEN_9716 = _T_3 ? _matrix_c_6_T_16 : _GEN_9701; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 296:24 327:27]
  wire [255:0] _GEN_9733 = _T_2 ? _GEN_9684 : _GEN_9706; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 296:24]
  wire [255:0] _GEN_9738 = _T_2 ? _GEN_9685 : _GEN_9711; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 296:24]
  wire [255:0] _GEN_9743 = _T_2 ? _GEN_9686 : _GEN_9716; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 296:24]
  wire [255:0] _GEN_9786 = _T_1 ? _GEN_9673 : _GEN_9733; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 296:24]
  wire [255:0] _GEN_9791 = _T_1 ? _GEN_9678 : _GEN_9738; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 296:24]
  wire [255:0] _GEN_9796 = _T_1 ? _GEN_9679 : _GEN_9743; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 296:24]
  wire [63:0] a_tile_v_162_1 = rf_a_tile_v_1_MPORT_162_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] a_tile_v_162_0 = rf_a_tile_v_0_MPORT_162_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_a_6_T_12 = {a_tile_v_162_1,a_tile_v_162_0,128'h0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 342:35]
  wire [63:0] matrix_b_6_tile_v_18_3 = rf_matrix_b_6_tile_v_3_MPORT_18_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_6_tile_v_18_2 = rf_matrix_b_6_tile_v_2_MPORT_18_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_6_tile_v_18_1 = rf_matrix_b_6_tile_v_1_MPORT_18_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_6_tile_v_18_0 = rf_matrix_b_6_tile_v_0_MPORT_18_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_b_6_T_18 = {matrix_b_6_tile_v_18_3,matrix_b_6_tile_v_18_2,matrix_b_6_tile_v_18_1,
    matrix_b_6_tile_v_18_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] matrix_c_6_tile_v_18_3 = rf_matrix_c_6_tile_v_3_MPORT_18_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_6_tile_v_18_2 = rf_matrix_c_6_tile_v_2_MPORT_18_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_6_tile_v_18_1 = rf_matrix_c_6_tile_v_1_MPORT_18_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_6_tile_v_18_0 = rf_matrix_c_6_tile_v_0_MPORT_18_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_c_6_T_18 = {matrix_c_6_tile_v_18_3,matrix_c_6_tile_v_18_2,matrix_c_6_tile_v_18_1,
    matrix_c_6_tile_v_18_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] a_tile_v_163_3 = rf_a_tile_v_3_MPORT_54_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] a_tile_v_163_2 = rf_a_tile_v_2_MPORT_54_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] a_tile_v_163_1 = rf_a_tile_v_1_MPORT_163_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] a_tile_v_163_0 = rf_a_tile_v_0_MPORT_163_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] a_163 = {a_tile_v_163_3,a_tile_v_163_2,a_tile_v_163_1,a_tile_v_163_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] matrix_b_6_tile_v_19_3 = rf_matrix_b_6_tile_v_3_MPORT_19_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_6_tile_v_19_2 = rf_matrix_b_6_tile_v_2_MPORT_19_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_6_tile_v_19_1 = rf_matrix_b_6_tile_v_1_MPORT_19_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_6_tile_v_19_0 = rf_matrix_b_6_tile_v_0_MPORT_19_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_b_6_T_19 = {matrix_b_6_tile_v_19_3,matrix_b_6_tile_v_19_2,matrix_b_6_tile_v_19_1,
    matrix_b_6_tile_v_19_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] matrix_c_6_tile_v_19_3 = rf_matrix_c_6_tile_v_3_MPORT_19_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_6_tile_v_19_2 = rf_matrix_c_6_tile_v_2_MPORT_19_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_6_tile_v_19_1 = rf_matrix_c_6_tile_v_1_MPORT_19_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_6_tile_v_19_0 = rf_matrix_c_6_tile_v_0_MPORT_19_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_c_6_T_19 = {matrix_c_6_tile_v_19_3,matrix_c_6_tile_v_19_2,matrix_c_6_tile_v_19_1,
    matrix_c_6_tile_v_19_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [255:0] _GEN_9861 = io_mixPc ? _matrix_a_6_T_12 : a_163; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 340:30 342:29 347:29]
  wire [255:0] _GEN_9866 = io_mixPc ? _matrix_b_6_T_18 : _matrix_b_6_T_19; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 340:30 343:29 348:29]
  wire [255:0] _GEN_9867 = io_mixPc ? _matrix_c_6_T_18 : _matrix_c_6_T_19; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 340:30 344:29 349:29]
  wire [63:0] a_tile_v_164_1 = rf_a_tile_v_1_MPORT_164_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] a_tile_v_164_0 = rf_a_tile_v_0_MPORT_164_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_a_6_T_13 = {a_tile_v_164_1,a_tile_v_164_0,128'h0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 355:35]
  wire [63:0] matrix_b_6_tile_v_20_3 = rf_matrix_b_6_tile_v_3_MPORT_20_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_6_tile_v_20_2 = rf_matrix_b_6_tile_v_2_MPORT_20_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_6_tile_v_20_1 = rf_matrix_b_6_tile_v_1_MPORT_20_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_6_tile_v_20_0 = rf_matrix_b_6_tile_v_0_MPORT_20_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_b_6_T_20 = {matrix_b_6_tile_v_20_3,matrix_b_6_tile_v_20_2,matrix_b_6_tile_v_20_1,
    matrix_b_6_tile_v_20_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] matrix_c_6_tile_v_20_3 = rf_matrix_c_6_tile_v_3_MPORT_20_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_6_tile_v_20_2 = rf_matrix_c_6_tile_v_2_MPORT_20_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_6_tile_v_20_1 = rf_matrix_c_6_tile_v_1_MPORT_20_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_6_tile_v_20_0 = rf_matrix_c_6_tile_v_0_MPORT_20_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_c_6_T_20 = {matrix_c_6_tile_v_20_3,matrix_c_6_tile_v_20_2,matrix_c_6_tile_v_20_1,
    matrix_c_6_tile_v_20_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] a_tile_v_165_3 = rf_a_tile_v_3_MPORT_55_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] a_tile_v_165_2 = rf_a_tile_v_2_MPORT_55_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] a_tile_v_165_1 = rf_a_tile_v_1_MPORT_165_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] a_tile_v_165_0 = rf_a_tile_v_0_MPORT_165_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] a_165 = {a_tile_v_165_3,a_tile_v_165_2,a_tile_v_165_1,a_tile_v_165_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] matrix_b_6_tile_v_21_3 = rf_matrix_b_6_tile_v_3_MPORT_21_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_6_tile_v_21_2 = rf_matrix_b_6_tile_v_2_MPORT_21_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_6_tile_v_21_1 = rf_matrix_b_6_tile_v_1_MPORT_21_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_6_tile_v_21_0 = rf_matrix_b_6_tile_v_0_MPORT_21_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_b_6_T_21 = {matrix_b_6_tile_v_21_3,matrix_b_6_tile_v_21_2,matrix_b_6_tile_v_21_1,
    matrix_b_6_tile_v_21_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] matrix_c_6_tile_v_21_3 = rf_matrix_c_6_tile_v_3_MPORT_21_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_6_tile_v_21_2 = rf_matrix_c_6_tile_v_2_MPORT_21_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_6_tile_v_21_1 = rf_matrix_c_6_tile_v_1_MPORT_21_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_6_tile_v_21_0 = rf_matrix_c_6_tile_v_0_MPORT_21_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_c_6_T_21 = {matrix_c_6_tile_v_21_3,matrix_c_6_tile_v_21_2,matrix_c_6_tile_v_21_1,
    matrix_c_6_tile_v_21_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [255:0] _GEN_9872 = io_mixPc ? _matrix_a_6_T_13 : a_165; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 353:30 355:29 360:29]
  wire [255:0] _GEN_9873 = io_mixPc ? _matrix_b_6_T_20 : _matrix_b_6_T_21; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 353:30 356:29 361:29]
  wire [255:0] _GEN_9874 = io_mixPc ? _matrix_c_6_T_20 : _matrix_c_6_T_21; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 353:30 357:29 362:29]
  wire [63:0] a_tile_v_166_1 = rf_a_tile_v_1_MPORT_166_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] a_tile_v_166_0 = rf_a_tile_v_0_MPORT_166_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_a_6_T_14 = {a_tile_v_166_1,a_tile_v_166_0,128'h0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 367:33]
  wire [63:0] matrix_b_6_tile_v_22_3 = rf_matrix_b_6_tile_v_3_MPORT_22_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_6_tile_v_22_2 = rf_matrix_b_6_tile_v_2_MPORT_22_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_6_tile_v_22_1 = rf_matrix_b_6_tile_v_1_MPORT_22_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_6_tile_v_22_0 = rf_matrix_b_6_tile_v_0_MPORT_22_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_b_6_T_22 = {matrix_b_6_tile_v_22_3,matrix_b_6_tile_v_22_2,matrix_b_6_tile_v_22_1,
    matrix_b_6_tile_v_22_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] matrix_c_6_tile_v_22_3 = rf_matrix_c_6_tile_v_3_MPORT_22_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_6_tile_v_22_2 = rf_matrix_c_6_tile_v_2_MPORT_22_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_6_tile_v_22_1 = rf_matrix_c_6_tile_v_1_MPORT_22_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_6_tile_v_22_0 = rf_matrix_c_6_tile_v_0_MPORT_22_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_c_6_T_22 = {matrix_c_6_tile_v_22_3,matrix_c_6_tile_v_22_2,matrix_c_6_tile_v_22_1,
    matrix_c_6_tile_v_22_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] a_tile_v_167_1 = rf_a_tile_v_1_MPORT_167_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] a_tile_v_167_0 = rf_a_tile_v_0_MPORT_167_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_a_6_T_15 = {a_tile_v_167_1,a_tile_v_167_0,128'h0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 373:33]
  wire [63:0] matrix_b_6_tile_v_23_3 = rf_matrix_b_6_tile_v_3_MPORT_23_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_6_tile_v_23_2 = rf_matrix_b_6_tile_v_2_MPORT_23_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_6_tile_v_23_1 = rf_matrix_b_6_tile_v_1_MPORT_23_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_6_tile_v_23_0 = rf_matrix_b_6_tile_v_0_MPORT_23_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_b_6_T_23 = {matrix_b_6_tile_v_23_3,matrix_b_6_tile_v_23_2,matrix_b_6_tile_v_23_1,
    matrix_b_6_tile_v_23_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] matrix_c_6_tile_v_23_3 = rf_matrix_c_6_tile_v_3_MPORT_23_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_6_tile_v_23_2 = rf_matrix_c_6_tile_v_2_MPORT_23_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_6_tile_v_23_1 = rf_matrix_c_6_tile_v_1_MPORT_23_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_6_tile_v_23_0 = rf_matrix_c_6_tile_v_0_MPORT_23_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_c_6_T_23 = {matrix_c_6_tile_v_23_3,matrix_c_6_tile_v_23_2,matrix_c_6_tile_v_23_1,
    matrix_c_6_tile_v_23_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [255:0] _GEN_9879 = _T_4 ? _matrix_a_6_T_15 : matrix_a_6; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 159:21 338:24 373:27]
  wire [255:0] _GEN_9884 = _T_4 ? _matrix_b_6_T_23 : matrix_b_6; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 160:21 338:24 374:27]
  wire [255:0] _GEN_9889 = _T_4 ? _matrix_c_6_T_23 : matrix_c_6; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 161:21 338:24 375:27]
  wire [255:0] _GEN_9894 = _T_3 ? _matrix_a_6_T_14 : _GEN_9879; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 338:24 367:27]
  wire [255:0] _GEN_9899 = _T_3 ? _matrix_b_6_T_22 : _GEN_9884; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 338:24 368:27]
  wire [255:0] _GEN_9904 = _T_3 ? _matrix_c_6_T_22 : _GEN_9889; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 338:24 369:27]
  wire [255:0] _GEN_9921 = _T_2 ? _GEN_9872 : _GEN_9894; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 338:24]
  wire [255:0] _GEN_9926 = _T_2 ? _GEN_9873 : _GEN_9899; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 338:24]
  wire [255:0] _GEN_9931 = _T_2 ? _GEN_9874 : _GEN_9904; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 338:24]
  wire [255:0] _GEN_9974 = _T_1 ? _GEN_9861 : _GEN_9921; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 338:24]
  wire [255:0] _GEN_9979 = _T_1 ? _GEN_9866 : _GEN_9926; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 338:24]
  wire [255:0] _GEN_9984 = _T_1 ? _GEN_9867 : _GEN_9931; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 338:24]
  wire [255:0] _GEN_10053 = 2'h3 == set ? _GEN_9974 : matrix_a_6; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 210:18 159:21]
  wire [255:0] _GEN_10058 = 2'h3 == set ? _GEN_9979 : matrix_b_6; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 210:18 160:21]
  wire [255:0] _GEN_10063 = 2'h3 == set ? _GEN_9984 : matrix_c_6; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 210:18 161:21]
  wire [63:0] a_tile_v_168_1 = rf_a_tile_v_1_MPORT_168_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] a_tile_v_168_0 = rf_a_tile_v_0_MPORT_168_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_a_7_T = {a_tile_v_168_1,a_tile_v_168_0,128'h0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 216:35]
  wire [63:0] matrix_b_7_tile_v__3 = rf_matrix_b_7_tile_v_3_MPORT_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_7_tile_v__2 = rf_matrix_b_7_tile_v_2_MPORT_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_7_tile_v__1 = rf_matrix_b_7_tile_v_1_MPORT_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_7_tile_v__0 = rf_matrix_b_7_tile_v_0_MPORT_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_b_7_T = {matrix_b_7_tile_v__3,matrix_b_7_tile_v__2,matrix_b_7_tile_v__1,matrix_b_7_tile_v__0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] matrix_c_7_tile_v__3 = rf_matrix_c_7_tile_v_3_MPORT_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_7_tile_v__2 = rf_matrix_c_7_tile_v_2_MPORT_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_7_tile_v__1 = rf_matrix_c_7_tile_v_1_MPORT_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_7_tile_v__0 = rf_matrix_c_7_tile_v_0_MPORT_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_c_7_T = {matrix_c_7_tile_v__3,matrix_c_7_tile_v__2,matrix_c_7_tile_v__1,matrix_c_7_tile_v__0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] a_tile_v_169_3 = rf_a_tile_v_3_MPORT_56_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] a_tile_v_169_2 = rf_a_tile_v_2_MPORT_56_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] a_tile_v_169_1 = rf_a_tile_v_1_MPORT_169_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] a_tile_v_169_0 = rf_a_tile_v_0_MPORT_169_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] a_169 = {a_tile_v_169_3,a_tile_v_169_2,a_tile_v_169_1,a_tile_v_169_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] matrix_b_7_tile_v_1_3 = rf_matrix_b_7_tile_v_3_MPORT_1_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_7_tile_v_1_2 = rf_matrix_b_7_tile_v_2_MPORT_1_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_7_tile_v_1_1 = rf_matrix_b_7_tile_v_1_MPORT_1_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_7_tile_v_1_0 = rf_matrix_b_7_tile_v_0_MPORT_1_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_b_7_T_1 = {matrix_b_7_tile_v_1_3,matrix_b_7_tile_v_1_2,matrix_b_7_tile_v_1_1,
    matrix_b_7_tile_v_1_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] matrix_c_7_tile_v_1_3 = rf_matrix_c_7_tile_v_3_MPORT_1_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_7_tile_v_1_2 = rf_matrix_c_7_tile_v_2_MPORT_1_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_7_tile_v_1_1 = rf_matrix_c_7_tile_v_1_MPORT_1_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_7_tile_v_1_0 = rf_matrix_c_7_tile_v_0_MPORT_1_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_c_7_T_1 = {matrix_c_7_tile_v_1_3,matrix_c_7_tile_v_1_2,matrix_c_7_tile_v_1_1,
    matrix_c_7_tile_v_1_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] a_tile_v_170_1 = rf_a_tile_v_1_MPORT_170_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] a_tile_v_170_0 = rf_a_tile_v_0_MPORT_170_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_a_7_T_1 = {a_tile_v_170_1,a_tile_v_170_0,128'h0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 229:35]
  wire [63:0] matrix_b_7_tile_v_2_3 = rf_matrix_b_7_tile_v_3_MPORT_2_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_7_tile_v_2_2 = rf_matrix_b_7_tile_v_2_MPORT_2_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_7_tile_v_2_1 = rf_matrix_b_7_tile_v_1_MPORT_2_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_7_tile_v_2_0 = rf_matrix_b_7_tile_v_0_MPORT_2_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_b_7_T_2 = {matrix_b_7_tile_v_2_3,matrix_b_7_tile_v_2_2,matrix_b_7_tile_v_2_1,
    matrix_b_7_tile_v_2_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] matrix_c_7_tile_v_2_3 = rf_matrix_c_7_tile_v_3_MPORT_2_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_7_tile_v_2_2 = rf_matrix_c_7_tile_v_2_MPORT_2_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_7_tile_v_2_1 = rf_matrix_c_7_tile_v_1_MPORT_2_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_7_tile_v_2_0 = rf_matrix_c_7_tile_v_0_MPORT_2_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_c_7_T_2 = {matrix_c_7_tile_v_2_3,matrix_c_7_tile_v_2_2,matrix_c_7_tile_v_2_1,
    matrix_c_7_tile_v_2_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] a_tile_v_171_3 = rf_a_tile_v_3_MPORT_57_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] a_tile_v_171_2 = rf_a_tile_v_2_MPORT_57_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] a_tile_v_171_1 = rf_a_tile_v_1_MPORT_171_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] a_tile_v_171_0 = rf_a_tile_v_0_MPORT_171_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] a_171 = {a_tile_v_171_3,a_tile_v_171_2,a_tile_v_171_1,a_tile_v_171_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] matrix_b_7_tile_v_3_3 = rf_matrix_b_7_tile_v_3_MPORT_3_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_7_tile_v_3_2 = rf_matrix_b_7_tile_v_2_MPORT_3_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_7_tile_v_3_1 = rf_matrix_b_7_tile_v_1_MPORT_3_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_7_tile_v_3_0 = rf_matrix_b_7_tile_v_0_MPORT_3_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_b_7_T_3 = {matrix_b_7_tile_v_3_3,matrix_b_7_tile_v_3_2,matrix_b_7_tile_v_3_1,
    matrix_b_7_tile_v_3_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] matrix_c_7_tile_v_3_3 = rf_matrix_c_7_tile_v_3_MPORT_3_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_7_tile_v_3_2 = rf_matrix_c_7_tile_v_2_MPORT_3_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_7_tile_v_3_1 = rf_matrix_c_7_tile_v_1_MPORT_3_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_7_tile_v_3_0 = rf_matrix_c_7_tile_v_0_MPORT_3_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_c_7_T_3 = {matrix_c_7_tile_v_3_3,matrix_c_7_tile_v_3_2,matrix_c_7_tile_v_3_1,
    matrix_c_7_tile_v_3_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [255:0] _GEN_10832 = io_mixPc ? _matrix_a_7_T_1 : a_171; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 227:30 229:29 234:29]
  wire [255:0] _GEN_10833 = io_mixPc ? _matrix_b_7_T_2 : _matrix_b_7_T_3; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 227:30 230:29 235:29]
  wire [255:0] _GEN_10838 = io_mixPc ? _matrix_c_7_T_2 : _matrix_c_7_T_3; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 227:30 231:29 236:29]
  wire [63:0] a_tile_v_172_1 = rf_a_tile_v_1_MPORT_172_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] a_tile_v_172_0 = rf_a_tile_v_0_MPORT_172_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_a_7_T_2 = {a_tile_v_172_1,a_tile_v_172_0,128'h0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 241:33]
  wire [63:0] matrix_b_7_tile_v_4_3 = rf_matrix_b_7_tile_v_3_MPORT_4_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_7_tile_v_4_2 = rf_matrix_b_7_tile_v_2_MPORT_4_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_7_tile_v_4_1 = rf_matrix_b_7_tile_v_1_MPORT_4_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_7_tile_v_4_0 = rf_matrix_b_7_tile_v_0_MPORT_4_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_b_7_T_4 = {matrix_b_7_tile_v_4_3,matrix_b_7_tile_v_4_2,matrix_b_7_tile_v_4_1,
    matrix_b_7_tile_v_4_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] matrix_c_7_tile_v_4_3 = rf_matrix_c_7_tile_v_3_MPORT_4_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_7_tile_v_4_2 = rf_matrix_c_7_tile_v_2_MPORT_4_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_7_tile_v_4_1 = rf_matrix_c_7_tile_v_1_MPORT_4_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_7_tile_v_4_0 = rf_matrix_c_7_tile_v_0_MPORT_4_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_c_7_T_4 = {matrix_c_7_tile_v_4_3,matrix_c_7_tile_v_4_2,matrix_c_7_tile_v_4_1,
    matrix_c_7_tile_v_4_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] a_tile_v_173_1 = rf_a_tile_v_1_MPORT_173_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] a_tile_v_173_0 = rf_a_tile_v_0_MPORT_173_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_a_7_T_3 = {a_tile_v_173_1,a_tile_v_173_0,128'h0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 247:33]
  wire [63:0] matrix_b_7_tile_v_5_3 = rf_matrix_b_7_tile_v_3_MPORT_5_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_7_tile_v_5_2 = rf_matrix_b_7_tile_v_2_MPORT_5_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_7_tile_v_5_1 = rf_matrix_b_7_tile_v_1_MPORT_5_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_7_tile_v_5_0 = rf_matrix_b_7_tile_v_0_MPORT_5_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_b_7_T_5 = {matrix_b_7_tile_v_5_3,matrix_b_7_tile_v_5_2,matrix_b_7_tile_v_5_1,
    matrix_b_7_tile_v_5_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] matrix_c_7_tile_v_5_3 = rf_matrix_c_7_tile_v_3_MPORT_5_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_7_tile_v_5_2 = rf_matrix_c_7_tile_v_2_MPORT_5_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_7_tile_v_5_1 = rf_matrix_c_7_tile_v_1_MPORT_5_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_7_tile_v_5_0 = rf_matrix_c_7_tile_v_0_MPORT_5_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_c_7_T_5 = {matrix_c_7_tile_v_5_3,matrix_c_7_tile_v_5_2,matrix_c_7_tile_v_5_1,
    matrix_c_7_tile_v_5_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [255:0] _GEN_10847 = 2'h3 == step ? _matrix_a_7_T_3 : matrix_a_7; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 159:21 212:23 247:27]
  wire [255:0] _GEN_10852 = 2'h3 == step ? _matrix_b_7_T_5 : matrix_b_7; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 160:21 212:23 248:27]
  wire [255:0] _GEN_10857 = 2'h3 == step ? _matrix_c_7_T_5 : matrix_c_7; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 161:21 212:23 249:27]
  wire [255:0] _GEN_10862 = 2'h2 == step ? _matrix_a_7_T_2 : _GEN_10847; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 212:23 241:27]
  wire [255:0] _GEN_10867 = 2'h2 == step ? _matrix_b_7_T_4 : _GEN_10852; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 212:23 242:27]
  wire [255:0] _GEN_10872 = 2'h2 == step ? _matrix_c_7_T_4 : _GEN_10857; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 212:23 243:27]
  wire [63:0] a_tile_v_174_1 = rf_a_tile_v_1_MPORT_174_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] a_tile_v_174_0 = rf_a_tile_v_0_MPORT_174_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_a_7_T_4 = {a_tile_v_174_1,a_tile_v_174_0,128'h0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 258:35]
  wire [63:0] matrix_b_7_tile_v_6_3 = rf_matrix_b_7_tile_v_3_MPORT_6_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_7_tile_v_6_2 = rf_matrix_b_7_tile_v_2_MPORT_6_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_7_tile_v_6_1 = rf_matrix_b_7_tile_v_1_MPORT_6_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_7_tile_v_6_0 = rf_matrix_b_7_tile_v_0_MPORT_6_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_b_7_T_6 = {matrix_b_7_tile_v_6_3,matrix_b_7_tile_v_6_2,matrix_b_7_tile_v_6_1,
    matrix_b_7_tile_v_6_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] matrix_c_7_tile_v_6_3 = rf_matrix_c_7_tile_v_3_MPORT_6_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_7_tile_v_6_2 = rf_matrix_c_7_tile_v_2_MPORT_6_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_7_tile_v_6_1 = rf_matrix_c_7_tile_v_1_MPORT_6_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_7_tile_v_6_0 = rf_matrix_c_7_tile_v_0_MPORT_6_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_c_7_T_6 = {matrix_c_7_tile_v_6_3,matrix_c_7_tile_v_6_2,matrix_c_7_tile_v_6_1,
    matrix_c_7_tile_v_6_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] a_tile_v_175_3 = rf_a_tile_v_3_MPORT_58_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] a_tile_v_175_2 = rf_a_tile_v_2_MPORT_58_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] a_tile_v_175_1 = rf_a_tile_v_1_MPORT_175_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] a_tile_v_175_0 = rf_a_tile_v_0_MPORT_175_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] a_175 = {a_tile_v_175_3,a_tile_v_175_2,a_tile_v_175_1,a_tile_v_175_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] matrix_b_7_tile_v_7_3 = rf_matrix_b_7_tile_v_3_MPORT_7_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_7_tile_v_7_2 = rf_matrix_b_7_tile_v_2_MPORT_7_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_7_tile_v_7_1 = rf_matrix_b_7_tile_v_1_MPORT_7_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_7_tile_v_7_0 = rf_matrix_b_7_tile_v_0_MPORT_7_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_b_7_T_7 = {matrix_b_7_tile_v_7_3,matrix_b_7_tile_v_7_2,matrix_b_7_tile_v_7_1,
    matrix_b_7_tile_v_7_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] matrix_c_7_tile_v_7_3 = rf_matrix_c_7_tile_v_3_MPORT_7_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_7_tile_v_7_2 = rf_matrix_c_7_tile_v_2_MPORT_7_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_7_tile_v_7_1 = rf_matrix_c_7_tile_v_1_MPORT_7_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_7_tile_v_7_0 = rf_matrix_c_7_tile_v_0_MPORT_7_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_c_7_T_7 = {matrix_c_7_tile_v_7_3,matrix_c_7_tile_v_7_2,matrix_c_7_tile_v_7_1,
    matrix_c_7_tile_v_7_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [255:0] _GEN_11017 = io_mixPc ? _matrix_a_7_T_4 : a_175; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 256:30 258:29 263:29]
  wire [255:0] _GEN_11018 = io_mixPc ? _matrix_b_7_T_6 : _matrix_b_7_T_7; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 256:30 259:29 264:29]
  wire [255:0] _GEN_11019 = io_mixPc ? _matrix_c_7_T_6 : _matrix_c_7_T_7; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 256:30 260:29 265:29]
  wire [63:0] a_tile_v_176_1 = rf_a_tile_v_1_MPORT_176_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] a_tile_v_176_0 = rf_a_tile_v_0_MPORT_176_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_a_7_T_5 = {a_tile_v_176_1,a_tile_v_176_0,128'h0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 271:35]
  wire [63:0] matrix_b_7_tile_v_8_3 = rf_matrix_b_7_tile_v_3_MPORT_8_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_7_tile_v_8_2 = rf_matrix_b_7_tile_v_2_MPORT_8_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_7_tile_v_8_1 = rf_matrix_b_7_tile_v_1_MPORT_8_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_7_tile_v_8_0 = rf_matrix_b_7_tile_v_0_MPORT_8_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_b_7_T_8 = {matrix_b_7_tile_v_8_3,matrix_b_7_tile_v_8_2,matrix_b_7_tile_v_8_1,
    matrix_b_7_tile_v_8_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] matrix_c_7_tile_v_8_3 = rf_matrix_c_7_tile_v_3_MPORT_8_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_7_tile_v_8_2 = rf_matrix_c_7_tile_v_2_MPORT_8_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_7_tile_v_8_1 = rf_matrix_c_7_tile_v_1_MPORT_8_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_7_tile_v_8_0 = rf_matrix_c_7_tile_v_0_MPORT_8_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_c_7_T_8 = {matrix_c_7_tile_v_8_3,matrix_c_7_tile_v_8_2,matrix_c_7_tile_v_8_1,
    matrix_c_7_tile_v_8_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] a_tile_v_177_3 = rf_a_tile_v_3_MPORT_59_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] a_tile_v_177_2 = rf_a_tile_v_2_MPORT_59_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] a_tile_v_177_1 = rf_a_tile_v_1_MPORT_177_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] a_tile_v_177_0 = rf_a_tile_v_0_MPORT_177_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] a_177 = {a_tile_v_177_3,a_tile_v_177_2,a_tile_v_177_1,a_tile_v_177_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] matrix_b_7_tile_v_9_3 = rf_matrix_b_7_tile_v_3_MPORT_9_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_7_tile_v_9_2 = rf_matrix_b_7_tile_v_2_MPORT_9_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_7_tile_v_9_1 = rf_matrix_b_7_tile_v_1_MPORT_9_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_7_tile_v_9_0 = rf_matrix_b_7_tile_v_0_MPORT_9_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_b_7_T_9 = {matrix_b_7_tile_v_9_3,matrix_b_7_tile_v_9_2,matrix_b_7_tile_v_9_1,
    matrix_b_7_tile_v_9_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] matrix_c_7_tile_v_9_3 = rf_matrix_c_7_tile_v_3_MPORT_9_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_7_tile_v_9_2 = rf_matrix_c_7_tile_v_2_MPORT_9_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_7_tile_v_9_1 = rf_matrix_c_7_tile_v_1_MPORT_9_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_7_tile_v_9_0 = rf_matrix_c_7_tile_v_0_MPORT_9_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_c_7_T_9 = {matrix_c_7_tile_v_9_3,matrix_c_7_tile_v_9_2,matrix_c_7_tile_v_9_1,
    matrix_c_7_tile_v_9_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [255:0] _GEN_11020 = io_mixPc ? _matrix_a_7_T_5 : a_177; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 269:30 271:29 276:29]
  wire [255:0] _GEN_11021 = io_mixPc ? _matrix_b_7_T_8 : _matrix_b_7_T_9; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 269:30 272:29 277:29]
  wire [255:0] _GEN_11022 = io_mixPc ? _matrix_c_7_T_8 : _matrix_c_7_T_9; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 269:30 273:29 278:29]
  wire [63:0] a_tile_v_178_1 = rf_a_tile_v_1_MPORT_178_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] a_tile_v_178_0 = rf_a_tile_v_0_MPORT_178_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_a_7_T_6 = {a_tile_v_178_1,a_tile_v_178_0,128'h0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 283:33]
  wire [63:0] matrix_b_7_tile_v_10_3 = rf_matrix_b_7_tile_v_3_MPORT_10_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_7_tile_v_10_2 = rf_matrix_b_7_tile_v_2_MPORT_10_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_7_tile_v_10_1 = rf_matrix_b_7_tile_v_1_MPORT_10_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_7_tile_v_10_0 = rf_matrix_b_7_tile_v_0_MPORT_10_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_b_7_T_10 = {matrix_b_7_tile_v_10_3,matrix_b_7_tile_v_10_2,matrix_b_7_tile_v_10_1,
    matrix_b_7_tile_v_10_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] matrix_c_7_tile_v_10_3 = rf_matrix_c_7_tile_v_3_MPORT_10_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_7_tile_v_10_2 = rf_matrix_c_7_tile_v_2_MPORT_10_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_7_tile_v_10_1 = rf_matrix_c_7_tile_v_1_MPORT_10_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_7_tile_v_10_0 = rf_matrix_c_7_tile_v_0_MPORT_10_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_c_7_T_10 = {matrix_c_7_tile_v_10_3,matrix_c_7_tile_v_10_2,matrix_c_7_tile_v_10_1,
    matrix_c_7_tile_v_10_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] a_tile_v_179_1 = rf_a_tile_v_1_MPORT_179_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] a_tile_v_179_0 = rf_a_tile_v_0_MPORT_179_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_a_7_T_7 = {a_tile_v_179_1,a_tile_v_179_0,128'h0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 289:33]
  wire [63:0] matrix_b_7_tile_v_11_3 = rf_matrix_b_7_tile_v_3_MPORT_11_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_7_tile_v_11_2 = rf_matrix_b_7_tile_v_2_MPORT_11_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_7_tile_v_11_1 = rf_matrix_b_7_tile_v_1_MPORT_11_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_7_tile_v_11_0 = rf_matrix_b_7_tile_v_0_MPORT_11_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_b_7_T_11 = {matrix_b_7_tile_v_11_3,matrix_b_7_tile_v_11_2,matrix_b_7_tile_v_11_1,
    matrix_b_7_tile_v_11_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] matrix_c_7_tile_v_11_3 = rf_matrix_c_7_tile_v_3_MPORT_11_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_7_tile_v_11_2 = rf_matrix_c_7_tile_v_2_MPORT_11_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_7_tile_v_11_1 = rf_matrix_c_7_tile_v_1_MPORT_11_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_7_tile_v_11_0 = rf_matrix_c_7_tile_v_0_MPORT_11_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_c_7_T_11 = {matrix_c_7_tile_v_11_3,matrix_c_7_tile_v_11_2,matrix_c_7_tile_v_11_1,
    matrix_c_7_tile_v_11_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [255:0] _GEN_11027 = _T_4 ? _matrix_a_7_T_7 : matrix_a_7; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 159:21 254:24 289:27]
  wire [255:0] _GEN_11032 = _T_4 ? _matrix_b_7_T_11 : matrix_b_7; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 160:21 254:24 290:27]
  wire [255:0] _GEN_11037 = _T_4 ? _matrix_c_7_T_11 : matrix_c_7; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 161:21 254:24 291:27]
  wire [255:0] _GEN_11042 = _T_3 ? _matrix_a_7_T_6 : _GEN_11027; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 254:24 283:27]
  wire [255:0] _GEN_11047 = _T_3 ? _matrix_b_7_T_10 : _GEN_11032; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 254:24 284:27]
  wire [255:0] _GEN_11052 = _T_3 ? _matrix_c_7_T_10 : _GEN_11037; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 254:24 285:27]
  wire [255:0] _GEN_11069 = _T_2 ? _GEN_11020 : _GEN_11042; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 254:24]
  wire [255:0] _GEN_11074 = _T_2 ? _GEN_11021 : _GEN_11047; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 254:24]
  wire [255:0] _GEN_11079 = _T_2 ? _GEN_11022 : _GEN_11052; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 254:24]
  wire [63:0] a_tile_v_180_1 = rf_a_tile_v_1_MPORT_180_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] a_tile_v_180_0 = rf_a_tile_v_0_MPORT_180_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_a_7_T_8 = {a_tile_v_180_1,a_tile_v_180_0,128'h0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 300:35]
  wire [63:0] matrix_b_7_tile_v_12_3 = rf_matrix_b_7_tile_v_3_MPORT_12_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_7_tile_v_12_2 = rf_matrix_b_7_tile_v_2_MPORT_12_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_7_tile_v_12_1 = rf_matrix_b_7_tile_v_1_MPORT_12_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_7_tile_v_12_0 = rf_matrix_b_7_tile_v_0_MPORT_12_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_b_7_T_12 = {matrix_b_7_tile_v_12_3,matrix_b_7_tile_v_12_2,matrix_b_7_tile_v_12_1,
    matrix_b_7_tile_v_12_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] matrix_c_7_tile_v_12_3 = rf_matrix_c_7_tile_v_3_MPORT_12_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_7_tile_v_12_2 = rf_matrix_c_7_tile_v_2_MPORT_12_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_7_tile_v_12_1 = rf_matrix_c_7_tile_v_1_MPORT_12_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_7_tile_v_12_0 = rf_matrix_c_7_tile_v_0_MPORT_12_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_c_7_T_12 = {matrix_c_7_tile_v_12_3,matrix_c_7_tile_v_12_2,matrix_c_7_tile_v_12_1,
    matrix_c_7_tile_v_12_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] a_tile_v_181_3 = rf_a_tile_v_3_MPORT_60_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] a_tile_v_181_2 = rf_a_tile_v_2_MPORT_60_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] a_tile_v_181_1 = rf_a_tile_v_1_MPORT_181_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] a_tile_v_181_0 = rf_a_tile_v_0_MPORT_181_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] a_181 = {a_tile_v_181_3,a_tile_v_181_2,a_tile_v_181_1,a_tile_v_181_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] matrix_b_7_tile_v_13_3 = rf_matrix_b_7_tile_v_3_MPORT_13_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_7_tile_v_13_2 = rf_matrix_b_7_tile_v_2_MPORT_13_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_7_tile_v_13_1 = rf_matrix_b_7_tile_v_1_MPORT_13_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_7_tile_v_13_0 = rf_matrix_b_7_tile_v_0_MPORT_13_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_b_7_T_13 = {matrix_b_7_tile_v_13_3,matrix_b_7_tile_v_13_2,matrix_b_7_tile_v_13_1,
    matrix_b_7_tile_v_13_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] matrix_c_7_tile_v_13_3 = rf_matrix_c_7_tile_v_3_MPORT_13_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_7_tile_v_13_2 = rf_matrix_c_7_tile_v_2_MPORT_13_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_7_tile_v_13_1 = rf_matrix_c_7_tile_v_1_MPORT_13_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_7_tile_v_13_0 = rf_matrix_c_7_tile_v_0_MPORT_13_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_c_7_T_13 = {matrix_c_7_tile_v_13_3,matrix_c_7_tile_v_13_2,matrix_c_7_tile_v_13_1,
    matrix_c_7_tile_v_13_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [255:0] _GEN_11197 = io_mixPc ? _matrix_a_7_T_8 : a_181; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 298:30 300:29 305:29]
  wire [255:0] _GEN_11198 = io_mixPc ? _matrix_b_7_T_12 : _matrix_b_7_T_13; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 298:30 301:29 306:29]
  wire [255:0] _GEN_11199 = io_mixPc ? _matrix_c_7_T_12 : _matrix_c_7_T_13; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 298:30 302:29 307:29]
  wire [63:0] a_tile_v_182_1 = rf_a_tile_v_1_MPORT_182_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] a_tile_v_182_0 = rf_a_tile_v_0_MPORT_182_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_a_7_T_9 = {a_tile_v_182_1,a_tile_v_182_0,128'h0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 313:35]
  wire [63:0] matrix_b_7_tile_v_14_3 = rf_matrix_b_7_tile_v_3_MPORT_14_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_7_tile_v_14_2 = rf_matrix_b_7_tile_v_2_MPORT_14_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_7_tile_v_14_1 = rf_matrix_b_7_tile_v_1_MPORT_14_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_7_tile_v_14_0 = rf_matrix_b_7_tile_v_0_MPORT_14_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_b_7_T_14 = {matrix_b_7_tile_v_14_3,matrix_b_7_tile_v_14_2,matrix_b_7_tile_v_14_1,
    matrix_b_7_tile_v_14_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] matrix_c_7_tile_v_14_3 = rf_matrix_c_7_tile_v_3_MPORT_14_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_7_tile_v_14_2 = rf_matrix_c_7_tile_v_2_MPORT_14_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_7_tile_v_14_1 = rf_matrix_c_7_tile_v_1_MPORT_14_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_7_tile_v_14_0 = rf_matrix_c_7_tile_v_0_MPORT_14_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_c_7_T_14 = {matrix_c_7_tile_v_14_3,matrix_c_7_tile_v_14_2,matrix_c_7_tile_v_14_1,
    matrix_c_7_tile_v_14_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] a_tile_v_183_3 = rf_a_tile_v_3_MPORT_61_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] a_tile_v_183_2 = rf_a_tile_v_2_MPORT_61_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] a_tile_v_183_1 = rf_a_tile_v_1_MPORT_183_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] a_tile_v_183_0 = rf_a_tile_v_0_MPORT_183_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] a_183 = {a_tile_v_183_3,a_tile_v_183_2,a_tile_v_183_1,a_tile_v_183_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] matrix_b_7_tile_v_15_3 = rf_matrix_b_7_tile_v_3_MPORT_15_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_7_tile_v_15_2 = rf_matrix_b_7_tile_v_2_MPORT_15_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_7_tile_v_15_1 = rf_matrix_b_7_tile_v_1_MPORT_15_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_7_tile_v_15_0 = rf_matrix_b_7_tile_v_0_MPORT_15_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_b_7_T_15 = {matrix_b_7_tile_v_15_3,matrix_b_7_tile_v_15_2,matrix_b_7_tile_v_15_1,
    matrix_b_7_tile_v_15_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] matrix_c_7_tile_v_15_3 = rf_matrix_c_7_tile_v_3_MPORT_15_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_7_tile_v_15_2 = rf_matrix_c_7_tile_v_2_MPORT_15_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_7_tile_v_15_1 = rf_matrix_c_7_tile_v_1_MPORT_15_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_7_tile_v_15_0 = rf_matrix_c_7_tile_v_0_MPORT_15_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_c_7_T_15 = {matrix_c_7_tile_v_15_3,matrix_c_7_tile_v_15_2,matrix_c_7_tile_v_15_1,
    matrix_c_7_tile_v_15_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [255:0] _GEN_11200 = io_mixPc ? _matrix_a_7_T_9 : a_183; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 311:30 313:29 318:29]
  wire [255:0] _GEN_11201 = io_mixPc ? _matrix_b_7_T_14 : _matrix_b_7_T_15; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 311:30 314:29 319:29]
  wire [255:0] _GEN_11202 = io_mixPc ? _matrix_c_7_T_14 : _matrix_c_7_T_15; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 311:30 315:29 320:29]
  wire [63:0] a_tile_v_184_1 = rf_a_tile_v_1_MPORT_184_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] a_tile_v_184_0 = rf_a_tile_v_0_MPORT_184_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_a_7_T_10 = {a_tile_v_184_1,a_tile_v_184_0,128'h0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 325:33]
  wire [63:0] matrix_b_7_tile_v_16_3 = rf_matrix_b_7_tile_v_3_MPORT_16_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_7_tile_v_16_2 = rf_matrix_b_7_tile_v_2_MPORT_16_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_7_tile_v_16_1 = rf_matrix_b_7_tile_v_1_MPORT_16_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_7_tile_v_16_0 = rf_matrix_b_7_tile_v_0_MPORT_16_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_b_7_T_16 = {matrix_b_7_tile_v_16_3,matrix_b_7_tile_v_16_2,matrix_b_7_tile_v_16_1,
    matrix_b_7_tile_v_16_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] matrix_c_7_tile_v_16_3 = rf_matrix_c_7_tile_v_3_MPORT_16_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_7_tile_v_16_2 = rf_matrix_c_7_tile_v_2_MPORT_16_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_7_tile_v_16_1 = rf_matrix_c_7_tile_v_1_MPORT_16_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_7_tile_v_16_0 = rf_matrix_c_7_tile_v_0_MPORT_16_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_c_7_T_16 = {matrix_c_7_tile_v_16_3,matrix_c_7_tile_v_16_2,matrix_c_7_tile_v_16_1,
    matrix_c_7_tile_v_16_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] a_tile_v_185_1 = rf_a_tile_v_1_MPORT_185_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] a_tile_v_185_0 = rf_a_tile_v_0_MPORT_185_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_a_7_T_11 = {a_tile_v_185_1,a_tile_v_185_0,128'h0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 331:33]
  wire [63:0] matrix_b_7_tile_v_17_3 = rf_matrix_b_7_tile_v_3_MPORT_17_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_7_tile_v_17_2 = rf_matrix_b_7_tile_v_2_MPORT_17_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_7_tile_v_17_1 = rf_matrix_b_7_tile_v_1_MPORT_17_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_7_tile_v_17_0 = rf_matrix_b_7_tile_v_0_MPORT_17_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_b_7_T_17 = {matrix_b_7_tile_v_17_3,matrix_b_7_tile_v_17_2,matrix_b_7_tile_v_17_1,
    matrix_b_7_tile_v_17_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] matrix_c_7_tile_v_17_3 = rf_matrix_c_7_tile_v_3_MPORT_17_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_7_tile_v_17_2 = rf_matrix_c_7_tile_v_2_MPORT_17_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_7_tile_v_17_1 = rf_matrix_c_7_tile_v_1_MPORT_17_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_7_tile_v_17_0 = rf_matrix_c_7_tile_v_0_MPORT_17_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_c_7_T_17 = {matrix_c_7_tile_v_17_3,matrix_c_7_tile_v_17_2,matrix_c_7_tile_v_17_1,
    matrix_c_7_tile_v_17_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [255:0] _GEN_11207 = _T_4 ? _matrix_a_7_T_11 : matrix_a_7; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 159:21 296:24 331:27]
  wire [255:0] _GEN_11212 = _T_4 ? _matrix_b_7_T_17 : matrix_b_7; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 160:21 296:24 332:27]
  wire [255:0] _GEN_11217 = _T_4 ? _matrix_c_7_T_17 : matrix_c_7; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 161:21 296:24 333:27]
  wire [255:0] _GEN_11222 = _T_3 ? _matrix_a_7_T_10 : _GEN_11207; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 296:24 325:27]
  wire [255:0] _GEN_11227 = _T_3 ? _matrix_b_7_T_16 : _GEN_11212; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 296:24 326:27]
  wire [255:0] _GEN_11232 = _T_3 ? _matrix_c_7_T_16 : _GEN_11217; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 296:24 327:27]
  wire [255:0] _GEN_11249 = _T_2 ? _GEN_11200 : _GEN_11222; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 296:24]
  wire [255:0] _GEN_11254 = _T_2 ? _GEN_11201 : _GEN_11227; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 296:24]
  wire [255:0] _GEN_11259 = _T_2 ? _GEN_11202 : _GEN_11232; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 296:24]
  wire [255:0] _GEN_11302 = _T_1 ? _GEN_11197 : _GEN_11249; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 296:24]
  wire [255:0] _GEN_11307 = _T_1 ? _GEN_11198 : _GEN_11254; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 296:24]
  wire [255:0] _GEN_11312 = _T_1 ? _GEN_11199 : _GEN_11259; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 296:24]
  wire [63:0] a_tile_v_186_1 = rf_a_tile_v_1_MPORT_186_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] a_tile_v_186_0 = rf_a_tile_v_0_MPORT_186_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_a_7_T_12 = {a_tile_v_186_1,a_tile_v_186_0,128'h0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 342:35]
  wire [63:0] matrix_b_7_tile_v_18_3 = rf_matrix_b_7_tile_v_3_MPORT_18_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_7_tile_v_18_2 = rf_matrix_b_7_tile_v_2_MPORT_18_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_7_tile_v_18_1 = rf_matrix_b_7_tile_v_1_MPORT_18_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_7_tile_v_18_0 = rf_matrix_b_7_tile_v_0_MPORT_18_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_b_7_T_18 = {matrix_b_7_tile_v_18_3,matrix_b_7_tile_v_18_2,matrix_b_7_tile_v_18_1,
    matrix_b_7_tile_v_18_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] matrix_c_7_tile_v_18_3 = rf_matrix_c_7_tile_v_3_MPORT_18_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_7_tile_v_18_2 = rf_matrix_c_7_tile_v_2_MPORT_18_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_7_tile_v_18_1 = rf_matrix_c_7_tile_v_1_MPORT_18_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_7_tile_v_18_0 = rf_matrix_c_7_tile_v_0_MPORT_18_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_c_7_T_18 = {matrix_c_7_tile_v_18_3,matrix_c_7_tile_v_18_2,matrix_c_7_tile_v_18_1,
    matrix_c_7_tile_v_18_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] a_tile_v_187_3 = rf_a_tile_v_3_MPORT_62_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] a_tile_v_187_2 = rf_a_tile_v_2_MPORT_62_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] a_tile_v_187_1 = rf_a_tile_v_1_MPORT_187_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] a_tile_v_187_0 = rf_a_tile_v_0_MPORT_187_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] a_187 = {a_tile_v_187_3,a_tile_v_187_2,a_tile_v_187_1,a_tile_v_187_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] matrix_b_7_tile_v_19_3 = rf_matrix_b_7_tile_v_3_MPORT_19_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_7_tile_v_19_2 = rf_matrix_b_7_tile_v_2_MPORT_19_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_7_tile_v_19_1 = rf_matrix_b_7_tile_v_1_MPORT_19_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_7_tile_v_19_0 = rf_matrix_b_7_tile_v_0_MPORT_19_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_b_7_T_19 = {matrix_b_7_tile_v_19_3,matrix_b_7_tile_v_19_2,matrix_b_7_tile_v_19_1,
    matrix_b_7_tile_v_19_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] matrix_c_7_tile_v_19_3 = rf_matrix_c_7_tile_v_3_MPORT_19_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_7_tile_v_19_2 = rf_matrix_c_7_tile_v_2_MPORT_19_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_7_tile_v_19_1 = rf_matrix_c_7_tile_v_1_MPORT_19_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_7_tile_v_19_0 = rf_matrix_c_7_tile_v_0_MPORT_19_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_c_7_T_19 = {matrix_c_7_tile_v_19_3,matrix_c_7_tile_v_19_2,matrix_c_7_tile_v_19_1,
    matrix_c_7_tile_v_19_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [255:0] _GEN_11377 = io_mixPc ? _matrix_a_7_T_12 : a_187; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 340:30 342:29 347:29]
  wire [255:0] _GEN_11378 = io_mixPc ? _matrix_b_7_T_18 : _matrix_b_7_T_19; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 340:30 343:29 348:29]
  wire [255:0] _GEN_11379 = io_mixPc ? _matrix_c_7_T_18 : _matrix_c_7_T_19; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 340:30 344:29 349:29]
  wire [63:0] a_tile_v_188_1 = rf_a_tile_v_1_MPORT_188_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] a_tile_v_188_0 = rf_a_tile_v_0_MPORT_188_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_a_7_T_13 = {a_tile_v_188_1,a_tile_v_188_0,128'h0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 355:35]
  wire [63:0] matrix_b_7_tile_v_20_3 = rf_matrix_b_7_tile_v_3_MPORT_20_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_7_tile_v_20_2 = rf_matrix_b_7_tile_v_2_MPORT_20_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_7_tile_v_20_1 = rf_matrix_b_7_tile_v_1_MPORT_20_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_7_tile_v_20_0 = rf_matrix_b_7_tile_v_0_MPORT_20_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_b_7_T_20 = {matrix_b_7_tile_v_20_3,matrix_b_7_tile_v_20_2,matrix_b_7_tile_v_20_1,
    matrix_b_7_tile_v_20_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] matrix_c_7_tile_v_20_3 = rf_matrix_c_7_tile_v_3_MPORT_20_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_7_tile_v_20_2 = rf_matrix_c_7_tile_v_2_MPORT_20_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_7_tile_v_20_1 = rf_matrix_c_7_tile_v_1_MPORT_20_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_7_tile_v_20_0 = rf_matrix_c_7_tile_v_0_MPORT_20_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_c_7_T_20 = {matrix_c_7_tile_v_20_3,matrix_c_7_tile_v_20_2,matrix_c_7_tile_v_20_1,
    matrix_c_7_tile_v_20_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] a_tile_v_189_3 = rf_a_tile_v_3_MPORT_63_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] a_tile_v_189_2 = rf_a_tile_v_2_MPORT_63_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] a_tile_v_189_1 = rf_a_tile_v_1_MPORT_189_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] a_tile_v_189_0 = rf_a_tile_v_0_MPORT_189_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] a_189 = {a_tile_v_189_3,a_tile_v_189_2,a_tile_v_189_1,a_tile_v_189_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] matrix_b_7_tile_v_21_3 = rf_matrix_b_7_tile_v_3_MPORT_21_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_7_tile_v_21_2 = rf_matrix_b_7_tile_v_2_MPORT_21_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_7_tile_v_21_1 = rf_matrix_b_7_tile_v_1_MPORT_21_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_7_tile_v_21_0 = rf_matrix_b_7_tile_v_0_MPORT_21_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_b_7_T_21 = {matrix_b_7_tile_v_21_3,matrix_b_7_tile_v_21_2,matrix_b_7_tile_v_21_1,
    matrix_b_7_tile_v_21_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] matrix_c_7_tile_v_21_3 = rf_matrix_c_7_tile_v_3_MPORT_21_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_7_tile_v_21_2 = rf_matrix_c_7_tile_v_2_MPORT_21_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_7_tile_v_21_1 = rf_matrix_c_7_tile_v_1_MPORT_21_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_7_tile_v_21_0 = rf_matrix_c_7_tile_v_0_MPORT_21_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_c_7_T_21 = {matrix_c_7_tile_v_21_3,matrix_c_7_tile_v_21_2,matrix_c_7_tile_v_21_1,
    matrix_c_7_tile_v_21_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [255:0] _GEN_11380 = io_mixPc ? _matrix_a_7_T_13 : a_189; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 353:30 355:29 360:29]
  wire [255:0] _GEN_11381 = io_mixPc ? _matrix_b_7_T_20 : _matrix_b_7_T_21; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 353:30 356:29 361:29]
  wire [255:0] _GEN_11382 = io_mixPc ? _matrix_c_7_T_20 : _matrix_c_7_T_21; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 353:30 357:29 362:29]
  wire [63:0] a_tile_v_190_1 = rf_a_tile_v_1_MPORT_190_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] a_tile_v_190_0 = rf_a_tile_v_0_MPORT_190_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_a_7_T_14 = {a_tile_v_190_1,a_tile_v_190_0,128'h0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 367:33]
  wire [63:0] matrix_b_7_tile_v_22_3 = rf_matrix_b_7_tile_v_3_MPORT_22_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_7_tile_v_22_2 = rf_matrix_b_7_tile_v_2_MPORT_22_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_7_tile_v_22_1 = rf_matrix_b_7_tile_v_1_MPORT_22_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_7_tile_v_22_0 = rf_matrix_b_7_tile_v_0_MPORT_22_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_b_7_T_22 = {matrix_b_7_tile_v_22_3,matrix_b_7_tile_v_22_2,matrix_b_7_tile_v_22_1,
    matrix_b_7_tile_v_22_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] matrix_c_7_tile_v_22_3 = rf_matrix_c_7_tile_v_3_MPORT_22_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_7_tile_v_22_2 = rf_matrix_c_7_tile_v_2_MPORT_22_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_7_tile_v_22_1 = rf_matrix_c_7_tile_v_1_MPORT_22_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_7_tile_v_22_0 = rf_matrix_c_7_tile_v_0_MPORT_22_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_c_7_T_22 = {matrix_c_7_tile_v_22_3,matrix_c_7_tile_v_22_2,matrix_c_7_tile_v_22_1,
    matrix_c_7_tile_v_22_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] a_tile_v_191_1 = rf_a_tile_v_1_MPORT_191_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] a_tile_v_191_0 = rf_a_tile_v_0_MPORT_191_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_a_7_T_15 = {a_tile_v_191_1,a_tile_v_191_0,128'h0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 373:33]
  wire [63:0] matrix_b_7_tile_v_23_3 = rf_matrix_b_7_tile_v_3_MPORT_23_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_7_tile_v_23_2 = rf_matrix_b_7_tile_v_2_MPORT_23_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_7_tile_v_23_1 = rf_matrix_b_7_tile_v_1_MPORT_23_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_b_7_tile_v_23_0 = rf_matrix_b_7_tile_v_0_MPORT_23_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_b_7_T_23 = {matrix_b_7_tile_v_23_3,matrix_b_7_tile_v_23_2,matrix_b_7_tile_v_23_1,
    matrix_b_7_tile_v_23_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [63:0] matrix_c_7_tile_v_23_3 = rf_matrix_c_7_tile_v_3_MPORT_23_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_7_tile_v_23_2 = rf_matrix_c_7_tile_v_2_MPORT_23_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_7_tile_v_23_1 = rf_matrix_c_7_tile_v_1_MPORT_23_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [63:0] matrix_c_7_tile_v_23_0 = rf_matrix_c_7_tile_v_0_MPORT_23_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  wire [255:0] _matrix_c_7_T_23 = {matrix_c_7_tile_v_23_3,matrix_c_7_tile_v_23_2,matrix_c_7_tile_v_23_1,
    matrix_c_7_tile_v_23_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 86:12]
  wire [255:0] _GEN_11387 = _T_4 ? _matrix_a_7_T_15 : matrix_a_7; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 159:21 338:24 373:27]
  wire [255:0] _GEN_11392 = _T_4 ? _matrix_b_7_T_23 : matrix_b_7; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 160:21 338:24 374:27]
  wire [255:0] _GEN_11397 = _T_4 ? _matrix_c_7_T_23 : matrix_c_7; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 161:21 338:24 375:27]
  wire [255:0] _GEN_11402 = _T_3 ? _matrix_a_7_T_14 : _GEN_11387; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 338:24 367:27]
  wire [255:0] _GEN_11407 = _T_3 ? _matrix_b_7_T_22 : _GEN_11392; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 338:24 368:27]
  wire [255:0] _GEN_11412 = _T_3 ? _matrix_c_7_T_22 : _GEN_11397; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 338:24 369:27]
  wire [255:0] _GEN_11429 = _T_2 ? _GEN_11380 : _GEN_11402; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 338:24]
  wire [255:0] _GEN_11434 = _T_2 ? _GEN_11381 : _GEN_11407; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 338:24]
  wire [255:0] _GEN_11439 = _T_2 ? _GEN_11382 : _GEN_11412; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 338:24]
  wire [255:0] _GEN_11482 = _T_1 ? _GEN_11377 : _GEN_11429; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 338:24]
  wire [255:0] _GEN_11487 = _T_1 ? _GEN_11378 : _GEN_11434; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 338:24]
  wire [255:0] _GEN_11492 = _T_1 ? _GEN_11379 : _GEN_11439; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 338:24]
  wire [255:0] _GEN_11561 = 2'h3 == set ? _GEN_11482 : matrix_a_7; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 210:18 159:21]
  wire [255:0] _GEN_11566 = 2'h3 == set ? _GEN_11487 : matrix_b_7; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 210:18 160:21]
  wire [255:0] _GEN_11571 = 2'h3 == set ? _GEN_11492 : matrix_c_7; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 210:18 161:21]
  wire [1:0] _set_T_1 = set + 2'h1; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 387:18]
  wire [1:0] _step_T_1 = step + 2'h1; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 389:20]
  wire  _T_162 = io_top_wb_ready & io_top_wb_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 52:35]
  wire  _GEN_15056 = 2'h2 == out_step ? 1'h0 : 2'h3 == out_step; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 394:21 8:15]
  wire  _GEN_15257 = 2'h1 == out_step ? 1'h0 : 2'h2 == out_step; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 394:21 8:15]
  wire  _GEN_15324 = 2'h1 == out_step ? 1'h0 : _GEN_15056; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 394:21 8:15]
  wire  _GEN_15391 = 2'h0 == out_step & io_mixPc; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 394:21 8:15]
  wire  _GEN_15458 = 2'h0 == out_step & _GEN_22; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 394:21 8:15]
  wire  _GEN_15525 = 2'h0 == out_step ? 1'h0 : 2'h1 == out_step & io_mixPc; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 394:21 8:15]
  wire  _GEN_15592 = 2'h0 == out_step ? 1'h0 : 2'h1 == out_step & _GEN_22; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 394:21 8:15]
  wire  _GEN_15659 = 2'h0 == out_step ? 1'h0 : _GEN_15257; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 394:21 8:15]
  wire  _GEN_15726 = 2'h0 == out_step ? 1'h0 : _GEN_15324; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 394:21 8:15]
  wire  _GEN_15791 = out_set == 2'h3 | _GEN_1; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 461:40 462:15]
  wire [1:0] _out_set_T_1 = out_set + 2'h1; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 464:26]
  wire [1:0] _out_step_T_1 = out_step + 2'h1; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 466:28]
  assign rf_a_tile_v_1_MPORT_en = handshaked & _GEN_1276;
  assign rf_a_tile_v_1_MPORT_addr = 8'h0;
  assign rf_a_tile_v_1_MPORT_data = rf[rf_a_tile_v_1_MPORT_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_0_MPORT_en = handshaked & _GEN_1276;
  assign rf_a_tile_v_0_MPORT_addr = 8'h4;
  assign rf_a_tile_v_0_MPORT_data = rf[rf_a_tile_v_0_MPORT_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_0_tile_v_3_MPORT_en = handshaked & _GEN_1276;
  assign rf_matrix_b_0_tile_v_3_MPORT_addr = 8'h40;
  assign rf_matrix_b_0_tile_v_3_MPORT_data = rf[rf_matrix_b_0_tile_v_3_MPORT_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_0_tile_v_2_MPORT_en = handshaked & _GEN_1276;
  assign rf_matrix_b_0_tile_v_2_MPORT_addr = 8'h44;
  assign rf_matrix_b_0_tile_v_2_MPORT_data = rf[rf_matrix_b_0_tile_v_2_MPORT_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_0_tile_v_1_MPORT_en = handshaked & _GEN_1276;
  assign rf_matrix_b_0_tile_v_1_MPORT_addr = 8'h48;
  assign rf_matrix_b_0_tile_v_1_MPORT_data = rf[rf_matrix_b_0_tile_v_1_MPORT_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_0_tile_v_0_MPORT_en = handshaked & _GEN_1276;
  assign rf_matrix_b_0_tile_v_0_MPORT_addr = 8'h4c;
  assign rf_matrix_b_0_tile_v_0_MPORT_data = rf[rf_matrix_b_0_tile_v_0_MPORT_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_0_tile_v_3_MPORT_en = handshaked & _GEN_1276;
  assign rf_matrix_c_0_tile_v_3_MPORT_addr = 8'h80;
  assign rf_matrix_c_0_tile_v_3_MPORT_data = rf[rf_matrix_c_0_tile_v_3_MPORT_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_0_tile_v_2_MPORT_en = handshaked & _GEN_1276;
  assign rf_matrix_c_0_tile_v_2_MPORT_addr = 8'h81;
  assign rf_matrix_c_0_tile_v_2_MPORT_data = rf[rf_matrix_c_0_tile_v_2_MPORT_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_0_tile_v_1_MPORT_en = handshaked & _GEN_1276;
  assign rf_matrix_c_0_tile_v_1_MPORT_addr = 8'h88;
  assign rf_matrix_c_0_tile_v_1_MPORT_data = rf[rf_matrix_c_0_tile_v_1_MPORT_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_0_tile_v_0_MPORT_en = handshaked & _GEN_1276;
  assign rf_matrix_c_0_tile_v_0_MPORT_addr = 8'h89;
  assign rf_matrix_c_0_tile_v_0_MPORT_data = rf[rf_matrix_c_0_tile_v_0_MPORT_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_3_MPORT_en = handshaked & _GEN_1291;
  assign rf_a_tile_v_3_MPORT_addr = 8'h0;
  assign rf_a_tile_v_3_MPORT_data = rf[rf_a_tile_v_3_MPORT_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_2_MPORT_en = handshaked & _GEN_1291;
  assign rf_a_tile_v_2_MPORT_addr = 8'h4;
  assign rf_a_tile_v_2_MPORT_data = rf[rf_a_tile_v_2_MPORT_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_1_MPORT_1_en = handshaked & _GEN_1291;
  assign rf_a_tile_v_1_MPORT_1_addr = 8'h8;
  assign rf_a_tile_v_1_MPORT_1_data = rf[rf_a_tile_v_1_MPORT_1_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_0_MPORT_1_en = handshaked & _GEN_1291;
  assign rf_a_tile_v_0_MPORT_1_addr = 8'hc;
  assign rf_a_tile_v_0_MPORT_1_data = rf[rf_a_tile_v_0_MPORT_1_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_0_tile_v_3_MPORT_1_en = handshaked & _GEN_1291;
  assign rf_matrix_b_0_tile_v_3_MPORT_1_addr = 8'h40;
  assign rf_matrix_b_0_tile_v_3_MPORT_1_data = rf[rf_matrix_b_0_tile_v_3_MPORT_1_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_0_tile_v_2_MPORT_1_en = handshaked & _GEN_1291;
  assign rf_matrix_b_0_tile_v_2_MPORT_1_addr = 8'h44;
  assign rf_matrix_b_0_tile_v_2_MPORT_1_data = rf[rf_matrix_b_0_tile_v_2_MPORT_1_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_0_tile_v_1_MPORT_1_en = handshaked & _GEN_1291;
  assign rf_matrix_b_0_tile_v_1_MPORT_1_addr = 8'h48;
  assign rf_matrix_b_0_tile_v_1_MPORT_1_data = rf[rf_matrix_b_0_tile_v_1_MPORT_1_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_0_tile_v_0_MPORT_1_en = handshaked & _GEN_1291;
  assign rf_matrix_b_0_tile_v_0_MPORT_1_addr = 8'h4c;
  assign rf_matrix_b_0_tile_v_0_MPORT_1_data = rf[rf_matrix_b_0_tile_v_0_MPORT_1_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_0_tile_v_3_MPORT_1_en = handshaked & _GEN_1291;
  assign rf_matrix_c_0_tile_v_3_MPORT_1_addr = 8'h80;
  assign rf_matrix_c_0_tile_v_3_MPORT_1_data = rf[rf_matrix_c_0_tile_v_3_MPORT_1_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_0_tile_v_2_MPORT_1_en = handshaked & _GEN_1291;
  assign rf_matrix_c_0_tile_v_2_MPORT_1_addr = 8'h84;
  assign rf_matrix_c_0_tile_v_2_MPORT_1_data = rf[rf_matrix_c_0_tile_v_2_MPORT_1_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_0_tile_v_1_MPORT_1_en = handshaked & _GEN_1291;
  assign rf_matrix_c_0_tile_v_1_MPORT_1_addr = 8'h88;
  assign rf_matrix_c_0_tile_v_1_MPORT_1_data = rf[rf_matrix_c_0_tile_v_1_MPORT_1_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_0_tile_v_0_MPORT_1_en = handshaked & _GEN_1291;
  assign rf_matrix_c_0_tile_v_0_MPORT_1_addr = 8'h8c;
  assign rf_matrix_c_0_tile_v_0_MPORT_1_data = rf[rf_matrix_c_0_tile_v_0_MPORT_1_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_1_MPORT_2_en = handshaked & _GEN_1305;
  assign rf_a_tile_v_1_MPORT_2_addr = 8'h8;
  assign rf_a_tile_v_1_MPORT_2_data = rf[rf_a_tile_v_1_MPORT_2_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_0_MPORT_2_en = handshaked & _GEN_1305;
  assign rf_a_tile_v_0_MPORT_2_addr = 8'hc;
  assign rf_a_tile_v_0_MPORT_2_data = rf[rf_a_tile_v_0_MPORT_2_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_0_tile_v_3_MPORT_2_en = handshaked & _GEN_1305;
  assign rf_matrix_b_0_tile_v_3_MPORT_2_addr = 8'h40;
  assign rf_matrix_b_0_tile_v_3_MPORT_2_data = rf[rf_matrix_b_0_tile_v_3_MPORT_2_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_0_tile_v_2_MPORT_2_en = handshaked & _GEN_1305;
  assign rf_matrix_b_0_tile_v_2_MPORT_2_addr = 8'h44;
  assign rf_matrix_b_0_tile_v_2_MPORT_2_data = rf[rf_matrix_b_0_tile_v_2_MPORT_2_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_0_tile_v_1_MPORT_2_en = handshaked & _GEN_1305;
  assign rf_matrix_b_0_tile_v_1_MPORT_2_addr = 8'h48;
  assign rf_matrix_b_0_tile_v_1_MPORT_2_data = rf[rf_matrix_b_0_tile_v_1_MPORT_2_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_0_tile_v_0_MPORT_2_en = handshaked & _GEN_1305;
  assign rf_matrix_b_0_tile_v_0_MPORT_2_addr = 8'h4c;
  assign rf_matrix_b_0_tile_v_0_MPORT_2_data = rf[rf_matrix_b_0_tile_v_0_MPORT_2_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_0_tile_v_3_MPORT_2_en = handshaked & _GEN_1305;
  assign rf_matrix_c_0_tile_v_3_MPORT_2_addr = 8'h90;
  assign rf_matrix_c_0_tile_v_3_MPORT_2_data = rf[rf_matrix_c_0_tile_v_3_MPORT_2_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_0_tile_v_2_MPORT_2_en = handshaked & _GEN_1305;
  assign rf_matrix_c_0_tile_v_2_MPORT_2_addr = 8'h91;
  assign rf_matrix_c_0_tile_v_2_MPORT_2_data = rf[rf_matrix_c_0_tile_v_2_MPORT_2_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_0_tile_v_1_MPORT_2_en = handshaked & _GEN_1305;
  assign rf_matrix_c_0_tile_v_1_MPORT_2_addr = 8'h98;
  assign rf_matrix_c_0_tile_v_1_MPORT_2_data = rf[rf_matrix_c_0_tile_v_1_MPORT_2_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_0_tile_v_0_MPORT_2_en = handshaked & _GEN_1305;
  assign rf_matrix_c_0_tile_v_0_MPORT_2_addr = 8'h99;
  assign rf_matrix_c_0_tile_v_0_MPORT_2_data = rf[rf_matrix_c_0_tile_v_0_MPORT_2_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_3_MPORT_1_en = handshaked & _GEN_1317;
  assign rf_a_tile_v_3_MPORT_1_addr = 8'h0;
  assign rf_a_tile_v_3_MPORT_1_data = rf[rf_a_tile_v_3_MPORT_1_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_2_MPORT_1_en = handshaked & _GEN_1317;
  assign rf_a_tile_v_2_MPORT_1_addr = 8'h4;
  assign rf_a_tile_v_2_MPORT_1_data = rf[rf_a_tile_v_2_MPORT_1_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_1_MPORT_3_en = handshaked & _GEN_1317;
  assign rf_a_tile_v_1_MPORT_3_addr = 8'h8;
  assign rf_a_tile_v_1_MPORT_3_data = rf[rf_a_tile_v_1_MPORT_3_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_0_MPORT_3_en = handshaked & _GEN_1317;
  assign rf_a_tile_v_0_MPORT_3_addr = 8'hc;
  assign rf_a_tile_v_0_MPORT_3_data = rf[rf_a_tile_v_0_MPORT_3_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_0_tile_v_3_MPORT_3_en = handshaked & _GEN_1317;
  assign rf_matrix_b_0_tile_v_3_MPORT_3_addr = 8'h40;
  assign rf_matrix_b_0_tile_v_3_MPORT_3_data = rf[rf_matrix_b_0_tile_v_3_MPORT_3_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_0_tile_v_2_MPORT_3_en = handshaked & _GEN_1317;
  assign rf_matrix_b_0_tile_v_2_MPORT_3_addr = 8'h44;
  assign rf_matrix_b_0_tile_v_2_MPORT_3_data = rf[rf_matrix_b_0_tile_v_2_MPORT_3_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_0_tile_v_1_MPORT_3_en = handshaked & _GEN_1317;
  assign rf_matrix_b_0_tile_v_1_MPORT_3_addr = 8'h48;
  assign rf_matrix_b_0_tile_v_1_MPORT_3_data = rf[rf_matrix_b_0_tile_v_1_MPORT_3_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_0_tile_v_0_MPORT_3_en = handshaked & _GEN_1317;
  assign rf_matrix_b_0_tile_v_0_MPORT_3_addr = 8'h4c;
  assign rf_matrix_b_0_tile_v_0_MPORT_3_data = rf[rf_matrix_b_0_tile_v_0_MPORT_3_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_0_tile_v_3_MPORT_3_en = handshaked & _GEN_1317;
  assign rf_matrix_c_0_tile_v_3_MPORT_3_addr = 8'h81;
  assign rf_matrix_c_0_tile_v_3_MPORT_3_data = rf[rf_matrix_c_0_tile_v_3_MPORT_3_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_0_tile_v_2_MPORT_3_en = handshaked & _GEN_1317;
  assign rf_matrix_c_0_tile_v_2_MPORT_3_addr = 8'h85;
  assign rf_matrix_c_0_tile_v_2_MPORT_3_data = rf[rf_matrix_c_0_tile_v_2_MPORT_3_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_0_tile_v_1_MPORT_3_en = handshaked & _GEN_1317;
  assign rf_matrix_c_0_tile_v_1_MPORT_3_addr = 8'h89;
  assign rf_matrix_c_0_tile_v_1_MPORT_3_data = rf[rf_matrix_c_0_tile_v_1_MPORT_3_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_0_tile_v_0_MPORT_3_en = handshaked & _GEN_1317;
  assign rf_matrix_c_0_tile_v_0_MPORT_3_addr = 8'h8d;
  assign rf_matrix_c_0_tile_v_0_MPORT_3_data = rf[rf_matrix_c_0_tile_v_0_MPORT_3_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_1_MPORT_4_en = handshaked & _GEN_1331;
  assign rf_a_tile_v_1_MPORT_4_addr = 8'h0;
  assign rf_a_tile_v_1_MPORT_4_data = rf[rf_a_tile_v_1_MPORT_4_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_0_MPORT_4_en = handshaked & _GEN_1331;
  assign rf_a_tile_v_0_MPORT_4_addr = 8'h4;
  assign rf_a_tile_v_0_MPORT_4_data = rf[rf_a_tile_v_0_MPORT_4_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_0_tile_v_3_MPORT_4_en = handshaked & _GEN_1331;
  assign rf_matrix_b_0_tile_v_3_MPORT_4_addr = 8'h40;
  assign rf_matrix_b_0_tile_v_3_MPORT_4_data = rf[rf_matrix_b_0_tile_v_3_MPORT_4_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_0_tile_v_2_MPORT_4_en = handshaked & _GEN_1331;
  assign rf_matrix_b_0_tile_v_2_MPORT_4_addr = 8'h44;
  assign rf_matrix_b_0_tile_v_2_MPORT_4_data = rf[rf_matrix_b_0_tile_v_2_MPORT_4_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_0_tile_v_1_MPORT_4_en = handshaked & _GEN_1331;
  assign rf_matrix_b_0_tile_v_1_MPORT_4_addr = 8'h48;
  assign rf_matrix_b_0_tile_v_1_MPORT_4_data = rf[rf_matrix_b_0_tile_v_1_MPORT_4_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_0_tile_v_0_MPORT_4_en = handshaked & _GEN_1331;
  assign rf_matrix_b_0_tile_v_0_MPORT_4_addr = 8'h4c;
  assign rf_matrix_b_0_tile_v_0_MPORT_4_data = rf[rf_matrix_b_0_tile_v_0_MPORT_4_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_0_tile_v_3_MPORT_4_en = handshaked & _GEN_1331;
  assign rf_matrix_c_0_tile_v_3_MPORT_4_addr = 8'h82;
  assign rf_matrix_c_0_tile_v_3_MPORT_4_data = rf[rf_matrix_c_0_tile_v_3_MPORT_4_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_0_tile_v_2_MPORT_4_en = handshaked & _GEN_1331;
  assign rf_matrix_c_0_tile_v_2_MPORT_4_addr = 8'h83;
  assign rf_matrix_c_0_tile_v_2_MPORT_4_data = rf[rf_matrix_c_0_tile_v_2_MPORT_4_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_0_tile_v_1_MPORT_4_en = handshaked & _GEN_1331;
  assign rf_matrix_c_0_tile_v_1_MPORT_4_addr = 8'h8a;
  assign rf_matrix_c_0_tile_v_1_MPORT_4_data = rf[rf_matrix_c_0_tile_v_1_MPORT_4_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_0_tile_v_0_MPORT_4_en = handshaked & _GEN_1331;
  assign rf_matrix_c_0_tile_v_0_MPORT_4_addr = 8'h8b;
  assign rf_matrix_c_0_tile_v_0_MPORT_4_data = rf[rf_matrix_c_0_tile_v_0_MPORT_4_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_1_MPORT_5_en = handshaked & _GEN_1343;
  assign rf_a_tile_v_1_MPORT_5_addr = 8'h8;
  assign rf_a_tile_v_1_MPORT_5_data = rf[rf_a_tile_v_1_MPORT_5_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_0_MPORT_5_en = handshaked & _GEN_1343;
  assign rf_a_tile_v_0_MPORT_5_addr = 8'hc;
  assign rf_a_tile_v_0_MPORT_5_data = rf[rf_a_tile_v_0_MPORT_5_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_0_tile_v_3_MPORT_5_en = handshaked & _GEN_1343;
  assign rf_matrix_b_0_tile_v_3_MPORT_5_addr = 8'h40;
  assign rf_matrix_b_0_tile_v_3_MPORT_5_data = rf[rf_matrix_b_0_tile_v_3_MPORT_5_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_0_tile_v_2_MPORT_5_en = handshaked & _GEN_1343;
  assign rf_matrix_b_0_tile_v_2_MPORT_5_addr = 8'h44;
  assign rf_matrix_b_0_tile_v_2_MPORT_5_data = rf[rf_matrix_b_0_tile_v_2_MPORT_5_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_0_tile_v_1_MPORT_5_en = handshaked & _GEN_1343;
  assign rf_matrix_b_0_tile_v_1_MPORT_5_addr = 8'h48;
  assign rf_matrix_b_0_tile_v_1_MPORT_5_data = rf[rf_matrix_b_0_tile_v_1_MPORT_5_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_0_tile_v_0_MPORT_5_en = handshaked & _GEN_1343;
  assign rf_matrix_b_0_tile_v_0_MPORT_5_addr = 8'h4c;
  assign rf_matrix_b_0_tile_v_0_MPORT_5_data = rf[rf_matrix_b_0_tile_v_0_MPORT_5_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_0_tile_v_3_MPORT_5_en = handshaked & _GEN_1343;
  assign rf_matrix_c_0_tile_v_3_MPORT_5_addr = 8'h92;
  assign rf_matrix_c_0_tile_v_3_MPORT_5_data = rf[rf_matrix_c_0_tile_v_3_MPORT_5_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_0_tile_v_2_MPORT_5_en = handshaked & _GEN_1343;
  assign rf_matrix_c_0_tile_v_2_MPORT_5_addr = 8'h93;
  assign rf_matrix_c_0_tile_v_2_MPORT_5_data = rf[rf_matrix_c_0_tile_v_2_MPORT_5_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_0_tile_v_1_MPORT_5_en = handshaked & _GEN_1343;
  assign rf_matrix_c_0_tile_v_1_MPORT_5_addr = 8'h9a;
  assign rf_matrix_c_0_tile_v_1_MPORT_5_data = rf[rf_matrix_c_0_tile_v_1_MPORT_5_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_0_tile_v_0_MPORT_5_en = handshaked & _GEN_1343;
  assign rf_matrix_c_0_tile_v_0_MPORT_5_addr = 8'h9b;
  assign rf_matrix_c_0_tile_v_0_MPORT_5_data = rf[rf_matrix_c_0_tile_v_0_MPORT_5_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_1_MPORT_6_en = handshaked & _GEN_1355;
  assign rf_a_tile_v_1_MPORT_6_addr = 8'h1;
  assign rf_a_tile_v_1_MPORT_6_data = rf[rf_a_tile_v_1_MPORT_6_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_0_MPORT_6_en = handshaked & _GEN_1355;
  assign rf_a_tile_v_0_MPORT_6_addr = 8'h5;
  assign rf_a_tile_v_0_MPORT_6_data = rf[rf_a_tile_v_0_MPORT_6_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_0_tile_v_3_MPORT_6_en = handshaked & _GEN_1355;
  assign rf_matrix_b_0_tile_v_3_MPORT_6_addr = 8'h50;
  assign rf_matrix_b_0_tile_v_3_MPORT_6_data = rf[rf_matrix_b_0_tile_v_3_MPORT_6_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_0_tile_v_2_MPORT_6_en = handshaked & _GEN_1355;
  assign rf_matrix_b_0_tile_v_2_MPORT_6_addr = 8'h54;
  assign rf_matrix_b_0_tile_v_2_MPORT_6_data = rf[rf_matrix_b_0_tile_v_2_MPORT_6_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_0_tile_v_1_MPORT_6_en = handshaked & _GEN_1355;
  assign rf_matrix_b_0_tile_v_1_MPORT_6_addr = 8'h58;
  assign rf_matrix_b_0_tile_v_1_MPORT_6_data = rf[rf_matrix_b_0_tile_v_1_MPORT_6_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_0_tile_v_0_MPORT_6_en = handshaked & _GEN_1355;
  assign rf_matrix_b_0_tile_v_0_MPORT_6_addr = 8'h5c;
  assign rf_matrix_b_0_tile_v_0_MPORT_6_data = rf[rf_matrix_b_0_tile_v_0_MPORT_6_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_0_tile_v_3_MPORT_6_en = handshaked & _GEN_1355;
  assign rf_matrix_c_0_tile_v_3_MPORT_6_addr = 8'h80;
  assign rf_matrix_c_0_tile_v_3_MPORT_6_data = rf[rf_matrix_c_0_tile_v_3_MPORT_6_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_0_tile_v_2_MPORT_6_en = handshaked & _GEN_1355;
  assign rf_matrix_c_0_tile_v_2_MPORT_6_addr = 8'h81;
  assign rf_matrix_c_0_tile_v_2_MPORT_6_data = rf[rf_matrix_c_0_tile_v_2_MPORT_6_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_0_tile_v_1_MPORT_6_en = handshaked & _GEN_1355;
  assign rf_matrix_c_0_tile_v_1_MPORT_6_addr = 8'h88;
  assign rf_matrix_c_0_tile_v_1_MPORT_6_data = rf[rf_matrix_c_0_tile_v_1_MPORT_6_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_0_tile_v_0_MPORT_6_en = handshaked & _GEN_1355;
  assign rf_matrix_c_0_tile_v_0_MPORT_6_addr = 8'h89;
  assign rf_matrix_c_0_tile_v_0_MPORT_6_data = rf[rf_matrix_c_0_tile_v_0_MPORT_6_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_3_MPORT_2_en = handshaked & _GEN_1367;
  assign rf_a_tile_v_3_MPORT_2_addr = 8'h1;
  assign rf_a_tile_v_3_MPORT_2_data = rf[rf_a_tile_v_3_MPORT_2_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_2_MPORT_2_en = handshaked & _GEN_1367;
  assign rf_a_tile_v_2_MPORT_2_addr = 8'h5;
  assign rf_a_tile_v_2_MPORT_2_data = rf[rf_a_tile_v_2_MPORT_2_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_1_MPORT_7_en = handshaked & _GEN_1367;
  assign rf_a_tile_v_1_MPORT_7_addr = 8'h9;
  assign rf_a_tile_v_1_MPORT_7_data = rf[rf_a_tile_v_1_MPORT_7_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_0_MPORT_7_en = handshaked & _GEN_1367;
  assign rf_a_tile_v_0_MPORT_7_addr = 8'hd;
  assign rf_a_tile_v_0_MPORT_7_data = rf[rf_a_tile_v_0_MPORT_7_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_0_tile_v_3_MPORT_7_en = handshaked & _GEN_1367;
  assign rf_matrix_b_0_tile_v_3_MPORT_7_addr = 8'h50;
  assign rf_matrix_b_0_tile_v_3_MPORT_7_data = rf[rf_matrix_b_0_tile_v_3_MPORT_7_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_0_tile_v_2_MPORT_7_en = handshaked & _GEN_1367;
  assign rf_matrix_b_0_tile_v_2_MPORT_7_addr = 8'h54;
  assign rf_matrix_b_0_tile_v_2_MPORT_7_data = rf[rf_matrix_b_0_tile_v_2_MPORT_7_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_0_tile_v_1_MPORT_7_en = handshaked & _GEN_1367;
  assign rf_matrix_b_0_tile_v_1_MPORT_7_addr = 8'h58;
  assign rf_matrix_b_0_tile_v_1_MPORT_7_data = rf[rf_matrix_b_0_tile_v_1_MPORT_7_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_0_tile_v_0_MPORT_7_en = handshaked & _GEN_1367;
  assign rf_matrix_b_0_tile_v_0_MPORT_7_addr = 8'h5c;
  assign rf_matrix_b_0_tile_v_0_MPORT_7_data = rf[rf_matrix_b_0_tile_v_0_MPORT_7_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_0_tile_v_3_MPORT_7_en = handshaked & _GEN_1367;
  assign rf_matrix_c_0_tile_v_3_MPORT_7_addr = 8'h80;
  assign rf_matrix_c_0_tile_v_3_MPORT_7_data = rf[rf_matrix_c_0_tile_v_3_MPORT_7_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_0_tile_v_2_MPORT_7_en = handshaked & _GEN_1367;
  assign rf_matrix_c_0_tile_v_2_MPORT_7_addr = 8'h84;
  assign rf_matrix_c_0_tile_v_2_MPORT_7_data = rf[rf_matrix_c_0_tile_v_2_MPORT_7_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_0_tile_v_1_MPORT_7_en = handshaked & _GEN_1367;
  assign rf_matrix_c_0_tile_v_1_MPORT_7_addr = 8'h88;
  assign rf_matrix_c_0_tile_v_1_MPORT_7_data = rf[rf_matrix_c_0_tile_v_1_MPORT_7_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_0_tile_v_0_MPORT_7_en = handshaked & _GEN_1367;
  assign rf_matrix_c_0_tile_v_0_MPORT_7_addr = 8'h8c;
  assign rf_matrix_c_0_tile_v_0_MPORT_7_data = rf[rf_matrix_c_0_tile_v_0_MPORT_7_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_1_MPORT_8_en = handshaked & _GEN_1381;
  assign rf_a_tile_v_1_MPORT_8_addr = 8'h9;
  assign rf_a_tile_v_1_MPORT_8_data = rf[rf_a_tile_v_1_MPORT_8_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_0_MPORT_8_en = handshaked & _GEN_1381;
  assign rf_a_tile_v_0_MPORT_8_addr = 8'hd;
  assign rf_a_tile_v_0_MPORT_8_data = rf[rf_a_tile_v_0_MPORT_8_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_0_tile_v_3_MPORT_8_en = handshaked & _GEN_1381;
  assign rf_matrix_b_0_tile_v_3_MPORT_8_addr = 8'h50;
  assign rf_matrix_b_0_tile_v_3_MPORT_8_data = rf[rf_matrix_b_0_tile_v_3_MPORT_8_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_0_tile_v_2_MPORT_8_en = handshaked & _GEN_1381;
  assign rf_matrix_b_0_tile_v_2_MPORT_8_addr = 8'h54;
  assign rf_matrix_b_0_tile_v_2_MPORT_8_data = rf[rf_matrix_b_0_tile_v_2_MPORT_8_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_0_tile_v_1_MPORT_8_en = handshaked & _GEN_1381;
  assign rf_matrix_b_0_tile_v_1_MPORT_8_addr = 8'h58;
  assign rf_matrix_b_0_tile_v_1_MPORT_8_data = rf[rf_matrix_b_0_tile_v_1_MPORT_8_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_0_tile_v_0_MPORT_8_en = handshaked & _GEN_1381;
  assign rf_matrix_b_0_tile_v_0_MPORT_8_addr = 8'h5c;
  assign rf_matrix_b_0_tile_v_0_MPORT_8_data = rf[rf_matrix_b_0_tile_v_0_MPORT_8_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_0_tile_v_3_MPORT_8_en = handshaked & _GEN_1381;
  assign rf_matrix_c_0_tile_v_3_MPORT_8_addr = 8'h90;
  assign rf_matrix_c_0_tile_v_3_MPORT_8_data = rf[rf_matrix_c_0_tile_v_3_MPORT_8_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_0_tile_v_2_MPORT_8_en = handshaked & _GEN_1381;
  assign rf_matrix_c_0_tile_v_2_MPORT_8_addr = 8'h91;
  assign rf_matrix_c_0_tile_v_2_MPORT_8_data = rf[rf_matrix_c_0_tile_v_2_MPORT_8_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_0_tile_v_1_MPORT_8_en = handshaked & _GEN_1381;
  assign rf_matrix_c_0_tile_v_1_MPORT_8_addr = 8'h98;
  assign rf_matrix_c_0_tile_v_1_MPORT_8_data = rf[rf_matrix_c_0_tile_v_1_MPORT_8_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_0_tile_v_0_MPORT_8_en = handshaked & _GEN_1381;
  assign rf_matrix_c_0_tile_v_0_MPORT_8_addr = 8'h99;
  assign rf_matrix_c_0_tile_v_0_MPORT_8_data = rf[rf_matrix_c_0_tile_v_0_MPORT_8_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_3_MPORT_3_en = handshaked & _GEN_1393;
  assign rf_a_tile_v_3_MPORT_3_addr = 8'h1;
  assign rf_a_tile_v_3_MPORT_3_data = rf[rf_a_tile_v_3_MPORT_3_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_2_MPORT_3_en = handshaked & _GEN_1393;
  assign rf_a_tile_v_2_MPORT_3_addr = 8'h5;
  assign rf_a_tile_v_2_MPORT_3_data = rf[rf_a_tile_v_2_MPORT_3_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_1_MPORT_9_en = handshaked & _GEN_1393;
  assign rf_a_tile_v_1_MPORT_9_addr = 8'h9;
  assign rf_a_tile_v_1_MPORT_9_data = rf[rf_a_tile_v_1_MPORT_9_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_0_MPORT_9_en = handshaked & _GEN_1393;
  assign rf_a_tile_v_0_MPORT_9_addr = 8'hd;
  assign rf_a_tile_v_0_MPORT_9_data = rf[rf_a_tile_v_0_MPORT_9_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_0_tile_v_3_MPORT_9_en = handshaked & _GEN_1393;
  assign rf_matrix_b_0_tile_v_3_MPORT_9_addr = 8'h50;
  assign rf_matrix_b_0_tile_v_3_MPORT_9_data = rf[rf_matrix_b_0_tile_v_3_MPORT_9_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_0_tile_v_2_MPORT_9_en = handshaked & _GEN_1393;
  assign rf_matrix_b_0_tile_v_2_MPORT_9_addr = 8'h54;
  assign rf_matrix_b_0_tile_v_2_MPORT_9_data = rf[rf_matrix_b_0_tile_v_2_MPORT_9_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_0_tile_v_1_MPORT_9_en = handshaked & _GEN_1393;
  assign rf_matrix_b_0_tile_v_1_MPORT_9_addr = 8'h58;
  assign rf_matrix_b_0_tile_v_1_MPORT_9_data = rf[rf_matrix_b_0_tile_v_1_MPORT_9_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_0_tile_v_0_MPORT_9_en = handshaked & _GEN_1393;
  assign rf_matrix_b_0_tile_v_0_MPORT_9_addr = 8'h5c;
  assign rf_matrix_b_0_tile_v_0_MPORT_9_data = rf[rf_matrix_b_0_tile_v_0_MPORT_9_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_0_tile_v_3_MPORT_9_en = handshaked & _GEN_1393;
  assign rf_matrix_c_0_tile_v_3_MPORT_9_addr = 8'h81;
  assign rf_matrix_c_0_tile_v_3_MPORT_9_data = rf[rf_matrix_c_0_tile_v_3_MPORT_9_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_0_tile_v_2_MPORT_9_en = handshaked & _GEN_1393;
  assign rf_matrix_c_0_tile_v_2_MPORT_9_addr = 8'h85;
  assign rf_matrix_c_0_tile_v_2_MPORT_9_data = rf[rf_matrix_c_0_tile_v_2_MPORT_9_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_0_tile_v_1_MPORT_9_en = handshaked & _GEN_1393;
  assign rf_matrix_c_0_tile_v_1_MPORT_9_addr = 8'h89;
  assign rf_matrix_c_0_tile_v_1_MPORT_9_data = rf[rf_matrix_c_0_tile_v_1_MPORT_9_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_0_tile_v_0_MPORT_9_en = handshaked & _GEN_1393;
  assign rf_matrix_c_0_tile_v_0_MPORT_9_addr = 8'h8d;
  assign rf_matrix_c_0_tile_v_0_MPORT_9_data = rf[rf_matrix_c_0_tile_v_0_MPORT_9_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_1_MPORT_10_en = handshaked & _GEN_1407;
  assign rf_a_tile_v_1_MPORT_10_addr = 8'h1;
  assign rf_a_tile_v_1_MPORT_10_data = rf[rf_a_tile_v_1_MPORT_10_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_0_MPORT_10_en = handshaked & _GEN_1407;
  assign rf_a_tile_v_0_MPORT_10_addr = 8'h5;
  assign rf_a_tile_v_0_MPORT_10_data = rf[rf_a_tile_v_0_MPORT_10_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_0_tile_v_3_MPORT_10_en = handshaked & _GEN_1407;
  assign rf_matrix_b_0_tile_v_3_MPORT_10_addr = 8'h50;
  assign rf_matrix_b_0_tile_v_3_MPORT_10_data = rf[rf_matrix_b_0_tile_v_3_MPORT_10_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_0_tile_v_2_MPORT_10_en = handshaked & _GEN_1407;
  assign rf_matrix_b_0_tile_v_2_MPORT_10_addr = 8'h54;
  assign rf_matrix_b_0_tile_v_2_MPORT_10_data = rf[rf_matrix_b_0_tile_v_2_MPORT_10_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_0_tile_v_1_MPORT_10_en = handshaked & _GEN_1407;
  assign rf_matrix_b_0_tile_v_1_MPORT_10_addr = 8'h58;
  assign rf_matrix_b_0_tile_v_1_MPORT_10_data = rf[rf_matrix_b_0_tile_v_1_MPORT_10_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_0_tile_v_0_MPORT_10_en = handshaked & _GEN_1407;
  assign rf_matrix_b_0_tile_v_0_MPORT_10_addr = 8'h5c;
  assign rf_matrix_b_0_tile_v_0_MPORT_10_data = rf[rf_matrix_b_0_tile_v_0_MPORT_10_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_0_tile_v_3_MPORT_10_en = handshaked & _GEN_1407;
  assign rf_matrix_c_0_tile_v_3_MPORT_10_addr = 8'h82;
  assign rf_matrix_c_0_tile_v_3_MPORT_10_data = rf[rf_matrix_c_0_tile_v_3_MPORT_10_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_0_tile_v_2_MPORT_10_en = handshaked & _GEN_1407;
  assign rf_matrix_c_0_tile_v_2_MPORT_10_addr = 8'h83;
  assign rf_matrix_c_0_tile_v_2_MPORT_10_data = rf[rf_matrix_c_0_tile_v_2_MPORT_10_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_0_tile_v_1_MPORT_10_en = handshaked & _GEN_1407;
  assign rf_matrix_c_0_tile_v_1_MPORT_10_addr = 8'h8a;
  assign rf_matrix_c_0_tile_v_1_MPORT_10_data = rf[rf_matrix_c_0_tile_v_1_MPORT_10_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_0_tile_v_0_MPORT_10_en = handshaked & _GEN_1407;
  assign rf_matrix_c_0_tile_v_0_MPORT_10_addr = 8'h8b;
  assign rf_matrix_c_0_tile_v_0_MPORT_10_data = rf[rf_matrix_c_0_tile_v_0_MPORT_10_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_1_MPORT_11_en = handshaked & _GEN_1419;
  assign rf_a_tile_v_1_MPORT_11_addr = 8'h9;
  assign rf_a_tile_v_1_MPORT_11_data = rf[rf_a_tile_v_1_MPORT_11_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_0_MPORT_11_en = handshaked & _GEN_1419;
  assign rf_a_tile_v_0_MPORT_11_addr = 8'hd;
  assign rf_a_tile_v_0_MPORT_11_data = rf[rf_a_tile_v_0_MPORT_11_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_0_tile_v_3_MPORT_11_en = handshaked & _GEN_1419;
  assign rf_matrix_b_0_tile_v_3_MPORT_11_addr = 8'h50;
  assign rf_matrix_b_0_tile_v_3_MPORT_11_data = rf[rf_matrix_b_0_tile_v_3_MPORT_11_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_0_tile_v_2_MPORT_11_en = handshaked & _GEN_1419;
  assign rf_matrix_b_0_tile_v_2_MPORT_11_addr = 8'h54;
  assign rf_matrix_b_0_tile_v_2_MPORT_11_data = rf[rf_matrix_b_0_tile_v_2_MPORT_11_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_0_tile_v_1_MPORT_11_en = handshaked & _GEN_1419;
  assign rf_matrix_b_0_tile_v_1_MPORT_11_addr = 8'h58;
  assign rf_matrix_b_0_tile_v_1_MPORT_11_data = rf[rf_matrix_b_0_tile_v_1_MPORT_11_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_0_tile_v_0_MPORT_11_en = handshaked & _GEN_1419;
  assign rf_matrix_b_0_tile_v_0_MPORT_11_addr = 8'h5c;
  assign rf_matrix_b_0_tile_v_0_MPORT_11_data = rf[rf_matrix_b_0_tile_v_0_MPORT_11_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_0_tile_v_3_MPORT_11_en = handshaked & _GEN_1419;
  assign rf_matrix_c_0_tile_v_3_MPORT_11_addr = 8'h92;
  assign rf_matrix_c_0_tile_v_3_MPORT_11_data = rf[rf_matrix_c_0_tile_v_3_MPORT_11_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_0_tile_v_2_MPORT_11_en = handshaked & _GEN_1419;
  assign rf_matrix_c_0_tile_v_2_MPORT_11_addr = 8'h93;
  assign rf_matrix_c_0_tile_v_2_MPORT_11_data = rf[rf_matrix_c_0_tile_v_2_MPORT_11_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_0_tile_v_1_MPORT_11_en = handshaked & _GEN_1419;
  assign rf_matrix_c_0_tile_v_1_MPORT_11_addr = 8'h9a;
  assign rf_matrix_c_0_tile_v_1_MPORT_11_data = rf[rf_matrix_c_0_tile_v_1_MPORT_11_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_0_tile_v_0_MPORT_11_en = handshaked & _GEN_1419;
  assign rf_matrix_c_0_tile_v_0_MPORT_11_addr = 8'h9b;
  assign rf_matrix_c_0_tile_v_0_MPORT_11_data = rf[rf_matrix_c_0_tile_v_0_MPORT_11_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_1_MPORT_12_en = handshaked & _GEN_1431;
  assign rf_a_tile_v_1_MPORT_12_addr = 8'h2;
  assign rf_a_tile_v_1_MPORT_12_data = rf[rf_a_tile_v_1_MPORT_12_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_0_MPORT_12_en = handshaked & _GEN_1431;
  assign rf_a_tile_v_0_MPORT_12_addr = 8'h6;
  assign rf_a_tile_v_0_MPORT_12_data = rf[rf_a_tile_v_0_MPORT_12_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_0_tile_v_3_MPORT_12_en = handshaked & _GEN_1431;
  assign rf_matrix_b_0_tile_v_3_MPORT_12_addr = 8'h60;
  assign rf_matrix_b_0_tile_v_3_MPORT_12_data = rf[rf_matrix_b_0_tile_v_3_MPORT_12_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_0_tile_v_2_MPORT_12_en = handshaked & _GEN_1431;
  assign rf_matrix_b_0_tile_v_2_MPORT_12_addr = 8'h64;
  assign rf_matrix_b_0_tile_v_2_MPORT_12_data = rf[rf_matrix_b_0_tile_v_2_MPORT_12_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_0_tile_v_1_MPORT_12_en = handshaked & _GEN_1431;
  assign rf_matrix_b_0_tile_v_1_MPORT_12_addr = 8'h68;
  assign rf_matrix_b_0_tile_v_1_MPORT_12_data = rf[rf_matrix_b_0_tile_v_1_MPORT_12_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_0_tile_v_0_MPORT_12_en = handshaked & _GEN_1431;
  assign rf_matrix_b_0_tile_v_0_MPORT_12_addr = 8'h6c;
  assign rf_matrix_b_0_tile_v_0_MPORT_12_data = rf[rf_matrix_b_0_tile_v_0_MPORT_12_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_0_tile_v_3_MPORT_12_en = handshaked & _GEN_1431;
  assign rf_matrix_c_0_tile_v_3_MPORT_12_addr = 8'h80;
  assign rf_matrix_c_0_tile_v_3_MPORT_12_data = rf[rf_matrix_c_0_tile_v_3_MPORT_12_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_0_tile_v_2_MPORT_12_en = handshaked & _GEN_1431;
  assign rf_matrix_c_0_tile_v_2_MPORT_12_addr = 8'h81;
  assign rf_matrix_c_0_tile_v_2_MPORT_12_data = rf[rf_matrix_c_0_tile_v_2_MPORT_12_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_0_tile_v_1_MPORT_12_en = handshaked & _GEN_1431;
  assign rf_matrix_c_0_tile_v_1_MPORT_12_addr = 8'h88;
  assign rf_matrix_c_0_tile_v_1_MPORT_12_data = rf[rf_matrix_c_0_tile_v_1_MPORT_12_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_0_tile_v_0_MPORT_12_en = handshaked & _GEN_1431;
  assign rf_matrix_c_0_tile_v_0_MPORT_12_addr = 8'h89;
  assign rf_matrix_c_0_tile_v_0_MPORT_12_data = rf[rf_matrix_c_0_tile_v_0_MPORT_12_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_3_MPORT_4_en = handshaked & _GEN_1443;
  assign rf_a_tile_v_3_MPORT_4_addr = 8'h2;
  assign rf_a_tile_v_3_MPORT_4_data = rf[rf_a_tile_v_3_MPORT_4_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_2_MPORT_4_en = handshaked & _GEN_1443;
  assign rf_a_tile_v_2_MPORT_4_addr = 8'h6;
  assign rf_a_tile_v_2_MPORT_4_data = rf[rf_a_tile_v_2_MPORT_4_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_1_MPORT_13_en = handshaked & _GEN_1443;
  assign rf_a_tile_v_1_MPORT_13_addr = 8'ha;
  assign rf_a_tile_v_1_MPORT_13_data = rf[rf_a_tile_v_1_MPORT_13_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_0_MPORT_13_en = handshaked & _GEN_1443;
  assign rf_a_tile_v_0_MPORT_13_addr = 8'he;
  assign rf_a_tile_v_0_MPORT_13_data = rf[rf_a_tile_v_0_MPORT_13_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_0_tile_v_3_MPORT_13_en = handshaked & _GEN_1443;
  assign rf_matrix_b_0_tile_v_3_MPORT_13_addr = 8'h60;
  assign rf_matrix_b_0_tile_v_3_MPORT_13_data = rf[rf_matrix_b_0_tile_v_3_MPORT_13_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_0_tile_v_2_MPORT_13_en = handshaked & _GEN_1443;
  assign rf_matrix_b_0_tile_v_2_MPORT_13_addr = 8'h64;
  assign rf_matrix_b_0_tile_v_2_MPORT_13_data = rf[rf_matrix_b_0_tile_v_2_MPORT_13_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_0_tile_v_1_MPORT_13_en = handshaked & _GEN_1443;
  assign rf_matrix_b_0_tile_v_1_MPORT_13_addr = 8'h68;
  assign rf_matrix_b_0_tile_v_1_MPORT_13_data = rf[rf_matrix_b_0_tile_v_1_MPORT_13_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_0_tile_v_0_MPORT_13_en = handshaked & _GEN_1443;
  assign rf_matrix_b_0_tile_v_0_MPORT_13_addr = 8'h6c;
  assign rf_matrix_b_0_tile_v_0_MPORT_13_data = rf[rf_matrix_b_0_tile_v_0_MPORT_13_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_0_tile_v_3_MPORT_13_en = handshaked & _GEN_1443;
  assign rf_matrix_c_0_tile_v_3_MPORT_13_addr = 8'h80;
  assign rf_matrix_c_0_tile_v_3_MPORT_13_data = rf[rf_matrix_c_0_tile_v_3_MPORT_13_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_0_tile_v_2_MPORT_13_en = handshaked & _GEN_1443;
  assign rf_matrix_c_0_tile_v_2_MPORT_13_addr = 8'h84;
  assign rf_matrix_c_0_tile_v_2_MPORT_13_data = rf[rf_matrix_c_0_tile_v_2_MPORT_13_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_0_tile_v_1_MPORT_13_en = handshaked & _GEN_1443;
  assign rf_matrix_c_0_tile_v_1_MPORT_13_addr = 8'h88;
  assign rf_matrix_c_0_tile_v_1_MPORT_13_data = rf[rf_matrix_c_0_tile_v_1_MPORT_13_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_0_tile_v_0_MPORT_13_en = handshaked & _GEN_1443;
  assign rf_matrix_c_0_tile_v_0_MPORT_13_addr = 8'h8c;
  assign rf_matrix_c_0_tile_v_0_MPORT_13_data = rf[rf_matrix_c_0_tile_v_0_MPORT_13_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_1_MPORT_14_en = handshaked & _GEN_1457;
  assign rf_a_tile_v_1_MPORT_14_addr = 8'ha;
  assign rf_a_tile_v_1_MPORT_14_data = rf[rf_a_tile_v_1_MPORT_14_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_0_MPORT_14_en = handshaked & _GEN_1457;
  assign rf_a_tile_v_0_MPORT_14_addr = 8'he;
  assign rf_a_tile_v_0_MPORT_14_data = rf[rf_a_tile_v_0_MPORT_14_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_0_tile_v_3_MPORT_14_en = handshaked & _GEN_1457;
  assign rf_matrix_b_0_tile_v_3_MPORT_14_addr = 8'h60;
  assign rf_matrix_b_0_tile_v_3_MPORT_14_data = rf[rf_matrix_b_0_tile_v_3_MPORT_14_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_0_tile_v_2_MPORT_14_en = handshaked & _GEN_1457;
  assign rf_matrix_b_0_tile_v_2_MPORT_14_addr = 8'h64;
  assign rf_matrix_b_0_tile_v_2_MPORT_14_data = rf[rf_matrix_b_0_tile_v_2_MPORT_14_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_0_tile_v_1_MPORT_14_en = handshaked & _GEN_1457;
  assign rf_matrix_b_0_tile_v_1_MPORT_14_addr = 8'h68;
  assign rf_matrix_b_0_tile_v_1_MPORT_14_data = rf[rf_matrix_b_0_tile_v_1_MPORT_14_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_0_tile_v_0_MPORT_14_en = handshaked & _GEN_1457;
  assign rf_matrix_b_0_tile_v_0_MPORT_14_addr = 8'h6c;
  assign rf_matrix_b_0_tile_v_0_MPORT_14_data = rf[rf_matrix_b_0_tile_v_0_MPORT_14_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_0_tile_v_3_MPORT_14_en = handshaked & _GEN_1457;
  assign rf_matrix_c_0_tile_v_3_MPORT_14_addr = 8'h90;
  assign rf_matrix_c_0_tile_v_3_MPORT_14_data = rf[rf_matrix_c_0_tile_v_3_MPORT_14_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_0_tile_v_2_MPORT_14_en = handshaked & _GEN_1457;
  assign rf_matrix_c_0_tile_v_2_MPORT_14_addr = 8'h91;
  assign rf_matrix_c_0_tile_v_2_MPORT_14_data = rf[rf_matrix_c_0_tile_v_2_MPORT_14_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_0_tile_v_1_MPORT_14_en = handshaked & _GEN_1457;
  assign rf_matrix_c_0_tile_v_1_MPORT_14_addr = 8'h98;
  assign rf_matrix_c_0_tile_v_1_MPORT_14_data = rf[rf_matrix_c_0_tile_v_1_MPORT_14_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_0_tile_v_0_MPORT_14_en = handshaked & _GEN_1457;
  assign rf_matrix_c_0_tile_v_0_MPORT_14_addr = 8'h99;
  assign rf_matrix_c_0_tile_v_0_MPORT_14_data = rf[rf_matrix_c_0_tile_v_0_MPORT_14_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_3_MPORT_5_en = handshaked & _GEN_1469;
  assign rf_a_tile_v_3_MPORT_5_addr = 8'h2;
  assign rf_a_tile_v_3_MPORT_5_data = rf[rf_a_tile_v_3_MPORT_5_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_2_MPORT_5_en = handshaked & _GEN_1469;
  assign rf_a_tile_v_2_MPORT_5_addr = 8'h6;
  assign rf_a_tile_v_2_MPORT_5_data = rf[rf_a_tile_v_2_MPORT_5_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_1_MPORT_15_en = handshaked & _GEN_1469;
  assign rf_a_tile_v_1_MPORT_15_addr = 8'ha;
  assign rf_a_tile_v_1_MPORT_15_data = rf[rf_a_tile_v_1_MPORT_15_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_0_MPORT_15_en = handshaked & _GEN_1469;
  assign rf_a_tile_v_0_MPORT_15_addr = 8'he;
  assign rf_a_tile_v_0_MPORT_15_data = rf[rf_a_tile_v_0_MPORT_15_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_0_tile_v_3_MPORT_15_en = handshaked & _GEN_1469;
  assign rf_matrix_b_0_tile_v_3_MPORT_15_addr = 8'h60;
  assign rf_matrix_b_0_tile_v_3_MPORT_15_data = rf[rf_matrix_b_0_tile_v_3_MPORT_15_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_0_tile_v_2_MPORT_15_en = handshaked & _GEN_1469;
  assign rf_matrix_b_0_tile_v_2_MPORT_15_addr = 8'h64;
  assign rf_matrix_b_0_tile_v_2_MPORT_15_data = rf[rf_matrix_b_0_tile_v_2_MPORT_15_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_0_tile_v_1_MPORT_15_en = handshaked & _GEN_1469;
  assign rf_matrix_b_0_tile_v_1_MPORT_15_addr = 8'h68;
  assign rf_matrix_b_0_tile_v_1_MPORT_15_data = rf[rf_matrix_b_0_tile_v_1_MPORT_15_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_0_tile_v_0_MPORT_15_en = handshaked & _GEN_1469;
  assign rf_matrix_b_0_tile_v_0_MPORT_15_addr = 8'h6c;
  assign rf_matrix_b_0_tile_v_0_MPORT_15_data = rf[rf_matrix_b_0_tile_v_0_MPORT_15_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_0_tile_v_3_MPORT_15_en = handshaked & _GEN_1469;
  assign rf_matrix_c_0_tile_v_3_MPORT_15_addr = 8'h81;
  assign rf_matrix_c_0_tile_v_3_MPORT_15_data = rf[rf_matrix_c_0_tile_v_3_MPORT_15_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_0_tile_v_2_MPORT_15_en = handshaked & _GEN_1469;
  assign rf_matrix_c_0_tile_v_2_MPORT_15_addr = 8'h85;
  assign rf_matrix_c_0_tile_v_2_MPORT_15_data = rf[rf_matrix_c_0_tile_v_2_MPORT_15_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_0_tile_v_1_MPORT_15_en = handshaked & _GEN_1469;
  assign rf_matrix_c_0_tile_v_1_MPORT_15_addr = 8'h89;
  assign rf_matrix_c_0_tile_v_1_MPORT_15_data = rf[rf_matrix_c_0_tile_v_1_MPORT_15_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_0_tile_v_0_MPORT_15_en = handshaked & _GEN_1469;
  assign rf_matrix_c_0_tile_v_0_MPORT_15_addr = 8'h8d;
  assign rf_matrix_c_0_tile_v_0_MPORT_15_data = rf[rf_matrix_c_0_tile_v_0_MPORT_15_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_1_MPORT_16_en = handshaked & _GEN_1483;
  assign rf_a_tile_v_1_MPORT_16_addr = 8'h2;
  assign rf_a_tile_v_1_MPORT_16_data = rf[rf_a_tile_v_1_MPORT_16_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_0_MPORT_16_en = handshaked & _GEN_1483;
  assign rf_a_tile_v_0_MPORT_16_addr = 8'h6;
  assign rf_a_tile_v_0_MPORT_16_data = rf[rf_a_tile_v_0_MPORT_16_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_0_tile_v_3_MPORT_16_en = handshaked & _GEN_1483;
  assign rf_matrix_b_0_tile_v_3_MPORT_16_addr = 8'h60;
  assign rf_matrix_b_0_tile_v_3_MPORT_16_data = rf[rf_matrix_b_0_tile_v_3_MPORT_16_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_0_tile_v_2_MPORT_16_en = handshaked & _GEN_1483;
  assign rf_matrix_b_0_tile_v_2_MPORT_16_addr = 8'h64;
  assign rf_matrix_b_0_tile_v_2_MPORT_16_data = rf[rf_matrix_b_0_tile_v_2_MPORT_16_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_0_tile_v_1_MPORT_16_en = handshaked & _GEN_1483;
  assign rf_matrix_b_0_tile_v_1_MPORT_16_addr = 8'h68;
  assign rf_matrix_b_0_tile_v_1_MPORT_16_data = rf[rf_matrix_b_0_tile_v_1_MPORT_16_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_0_tile_v_0_MPORT_16_en = handshaked & _GEN_1483;
  assign rf_matrix_b_0_tile_v_0_MPORT_16_addr = 8'h6c;
  assign rf_matrix_b_0_tile_v_0_MPORT_16_data = rf[rf_matrix_b_0_tile_v_0_MPORT_16_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_0_tile_v_3_MPORT_16_en = handshaked & _GEN_1483;
  assign rf_matrix_c_0_tile_v_3_MPORT_16_addr = 8'h82;
  assign rf_matrix_c_0_tile_v_3_MPORT_16_data = rf[rf_matrix_c_0_tile_v_3_MPORT_16_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_0_tile_v_2_MPORT_16_en = handshaked & _GEN_1483;
  assign rf_matrix_c_0_tile_v_2_MPORT_16_addr = 8'h83;
  assign rf_matrix_c_0_tile_v_2_MPORT_16_data = rf[rf_matrix_c_0_tile_v_2_MPORT_16_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_0_tile_v_1_MPORT_16_en = handshaked & _GEN_1483;
  assign rf_matrix_c_0_tile_v_1_MPORT_16_addr = 8'h8a;
  assign rf_matrix_c_0_tile_v_1_MPORT_16_data = rf[rf_matrix_c_0_tile_v_1_MPORT_16_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_0_tile_v_0_MPORT_16_en = handshaked & _GEN_1483;
  assign rf_matrix_c_0_tile_v_0_MPORT_16_addr = 8'h8b;
  assign rf_matrix_c_0_tile_v_0_MPORT_16_data = rf[rf_matrix_c_0_tile_v_0_MPORT_16_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_1_MPORT_17_en = handshaked & _GEN_1495;
  assign rf_a_tile_v_1_MPORT_17_addr = 8'ha;
  assign rf_a_tile_v_1_MPORT_17_data = rf[rf_a_tile_v_1_MPORT_17_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_0_MPORT_17_en = handshaked & _GEN_1495;
  assign rf_a_tile_v_0_MPORT_17_addr = 8'he;
  assign rf_a_tile_v_0_MPORT_17_data = rf[rf_a_tile_v_0_MPORT_17_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_0_tile_v_3_MPORT_17_en = handshaked & _GEN_1495;
  assign rf_matrix_b_0_tile_v_3_MPORT_17_addr = 8'h60;
  assign rf_matrix_b_0_tile_v_3_MPORT_17_data = rf[rf_matrix_b_0_tile_v_3_MPORT_17_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_0_tile_v_2_MPORT_17_en = handshaked & _GEN_1495;
  assign rf_matrix_b_0_tile_v_2_MPORT_17_addr = 8'h64;
  assign rf_matrix_b_0_tile_v_2_MPORT_17_data = rf[rf_matrix_b_0_tile_v_2_MPORT_17_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_0_tile_v_1_MPORT_17_en = handshaked & _GEN_1495;
  assign rf_matrix_b_0_tile_v_1_MPORT_17_addr = 8'h68;
  assign rf_matrix_b_0_tile_v_1_MPORT_17_data = rf[rf_matrix_b_0_tile_v_1_MPORT_17_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_0_tile_v_0_MPORT_17_en = handshaked & _GEN_1495;
  assign rf_matrix_b_0_tile_v_0_MPORT_17_addr = 8'h6c;
  assign rf_matrix_b_0_tile_v_0_MPORT_17_data = rf[rf_matrix_b_0_tile_v_0_MPORT_17_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_0_tile_v_3_MPORT_17_en = handshaked & _GEN_1495;
  assign rf_matrix_c_0_tile_v_3_MPORT_17_addr = 8'h92;
  assign rf_matrix_c_0_tile_v_3_MPORT_17_data = rf[rf_matrix_c_0_tile_v_3_MPORT_17_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_0_tile_v_2_MPORT_17_en = handshaked & _GEN_1495;
  assign rf_matrix_c_0_tile_v_2_MPORT_17_addr = 8'h93;
  assign rf_matrix_c_0_tile_v_2_MPORT_17_data = rf[rf_matrix_c_0_tile_v_2_MPORT_17_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_0_tile_v_1_MPORT_17_en = handshaked & _GEN_1495;
  assign rf_matrix_c_0_tile_v_1_MPORT_17_addr = 8'h9a;
  assign rf_matrix_c_0_tile_v_1_MPORT_17_data = rf[rf_matrix_c_0_tile_v_1_MPORT_17_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_0_tile_v_0_MPORT_17_en = handshaked & _GEN_1495;
  assign rf_matrix_c_0_tile_v_0_MPORT_17_addr = 8'h9b;
  assign rf_matrix_c_0_tile_v_0_MPORT_17_data = rf[rf_matrix_c_0_tile_v_0_MPORT_17_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_1_MPORT_18_en = handshaked & _GEN_1507;
  assign rf_a_tile_v_1_MPORT_18_addr = 8'h3;
  assign rf_a_tile_v_1_MPORT_18_data = rf[rf_a_tile_v_1_MPORT_18_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_0_MPORT_18_en = handshaked & _GEN_1507;
  assign rf_a_tile_v_0_MPORT_18_addr = 8'h7;
  assign rf_a_tile_v_0_MPORT_18_data = rf[rf_a_tile_v_0_MPORT_18_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_0_tile_v_3_MPORT_18_en = handshaked & _GEN_1507;
  assign rf_matrix_b_0_tile_v_3_MPORT_18_addr = 8'h70;
  assign rf_matrix_b_0_tile_v_3_MPORT_18_data = rf[rf_matrix_b_0_tile_v_3_MPORT_18_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_0_tile_v_2_MPORT_18_en = handshaked & _GEN_1507;
  assign rf_matrix_b_0_tile_v_2_MPORT_18_addr = 8'h74;
  assign rf_matrix_b_0_tile_v_2_MPORT_18_data = rf[rf_matrix_b_0_tile_v_2_MPORT_18_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_0_tile_v_1_MPORT_18_en = handshaked & _GEN_1507;
  assign rf_matrix_b_0_tile_v_1_MPORT_18_addr = 8'h78;
  assign rf_matrix_b_0_tile_v_1_MPORT_18_data = rf[rf_matrix_b_0_tile_v_1_MPORT_18_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_0_tile_v_0_MPORT_18_en = handshaked & _GEN_1507;
  assign rf_matrix_b_0_tile_v_0_MPORT_18_addr = 8'h7c;
  assign rf_matrix_b_0_tile_v_0_MPORT_18_data = rf[rf_matrix_b_0_tile_v_0_MPORT_18_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_0_tile_v_3_MPORT_18_en = handshaked & _GEN_1507;
  assign rf_matrix_c_0_tile_v_3_MPORT_18_addr = 8'h80;
  assign rf_matrix_c_0_tile_v_3_MPORT_18_data = rf[rf_matrix_c_0_tile_v_3_MPORT_18_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_0_tile_v_2_MPORT_18_en = handshaked & _GEN_1507;
  assign rf_matrix_c_0_tile_v_2_MPORT_18_addr = 8'h81;
  assign rf_matrix_c_0_tile_v_2_MPORT_18_data = rf[rf_matrix_c_0_tile_v_2_MPORT_18_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_0_tile_v_1_MPORT_18_en = handshaked & _GEN_1507;
  assign rf_matrix_c_0_tile_v_1_MPORT_18_addr = 8'h88;
  assign rf_matrix_c_0_tile_v_1_MPORT_18_data = rf[rf_matrix_c_0_tile_v_1_MPORT_18_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_0_tile_v_0_MPORT_18_en = handshaked & _GEN_1507;
  assign rf_matrix_c_0_tile_v_0_MPORT_18_addr = 8'h89;
  assign rf_matrix_c_0_tile_v_0_MPORT_18_data = rf[rf_matrix_c_0_tile_v_0_MPORT_18_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_3_MPORT_6_en = handshaked & _GEN_1519;
  assign rf_a_tile_v_3_MPORT_6_addr = 8'h3;
  assign rf_a_tile_v_3_MPORT_6_data = rf[rf_a_tile_v_3_MPORT_6_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_2_MPORT_6_en = handshaked & _GEN_1519;
  assign rf_a_tile_v_2_MPORT_6_addr = 8'h7;
  assign rf_a_tile_v_2_MPORT_6_data = rf[rf_a_tile_v_2_MPORT_6_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_1_MPORT_19_en = handshaked & _GEN_1519;
  assign rf_a_tile_v_1_MPORT_19_addr = 8'hb;
  assign rf_a_tile_v_1_MPORT_19_data = rf[rf_a_tile_v_1_MPORT_19_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_0_MPORT_19_en = handshaked & _GEN_1519;
  assign rf_a_tile_v_0_MPORT_19_addr = 8'hf;
  assign rf_a_tile_v_0_MPORT_19_data = rf[rf_a_tile_v_0_MPORT_19_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_0_tile_v_3_MPORT_19_en = handshaked & _GEN_1519;
  assign rf_matrix_b_0_tile_v_3_MPORT_19_addr = 8'h70;
  assign rf_matrix_b_0_tile_v_3_MPORT_19_data = rf[rf_matrix_b_0_tile_v_3_MPORT_19_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_0_tile_v_2_MPORT_19_en = handshaked & _GEN_1519;
  assign rf_matrix_b_0_tile_v_2_MPORT_19_addr = 8'h74;
  assign rf_matrix_b_0_tile_v_2_MPORT_19_data = rf[rf_matrix_b_0_tile_v_2_MPORT_19_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_0_tile_v_1_MPORT_19_en = handshaked & _GEN_1519;
  assign rf_matrix_b_0_tile_v_1_MPORT_19_addr = 8'h78;
  assign rf_matrix_b_0_tile_v_1_MPORT_19_data = rf[rf_matrix_b_0_tile_v_1_MPORT_19_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_0_tile_v_0_MPORT_19_en = handshaked & _GEN_1519;
  assign rf_matrix_b_0_tile_v_0_MPORT_19_addr = 8'h7c;
  assign rf_matrix_b_0_tile_v_0_MPORT_19_data = rf[rf_matrix_b_0_tile_v_0_MPORT_19_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_0_tile_v_3_MPORT_19_en = handshaked & _GEN_1519;
  assign rf_matrix_c_0_tile_v_3_MPORT_19_addr = 8'h80;
  assign rf_matrix_c_0_tile_v_3_MPORT_19_data = rf[rf_matrix_c_0_tile_v_3_MPORT_19_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_0_tile_v_2_MPORT_19_en = handshaked & _GEN_1519;
  assign rf_matrix_c_0_tile_v_2_MPORT_19_addr = 8'h84;
  assign rf_matrix_c_0_tile_v_2_MPORT_19_data = rf[rf_matrix_c_0_tile_v_2_MPORT_19_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_0_tile_v_1_MPORT_19_en = handshaked & _GEN_1519;
  assign rf_matrix_c_0_tile_v_1_MPORT_19_addr = 8'h88;
  assign rf_matrix_c_0_tile_v_1_MPORT_19_data = rf[rf_matrix_c_0_tile_v_1_MPORT_19_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_0_tile_v_0_MPORT_19_en = handshaked & _GEN_1519;
  assign rf_matrix_c_0_tile_v_0_MPORT_19_addr = 8'h8c;
  assign rf_matrix_c_0_tile_v_0_MPORT_19_data = rf[rf_matrix_c_0_tile_v_0_MPORT_19_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_1_MPORT_20_en = handshaked & _GEN_1533;
  assign rf_a_tile_v_1_MPORT_20_addr = 8'hb;
  assign rf_a_tile_v_1_MPORT_20_data = rf[rf_a_tile_v_1_MPORT_20_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_0_MPORT_20_en = handshaked & _GEN_1533;
  assign rf_a_tile_v_0_MPORT_20_addr = 8'hf;
  assign rf_a_tile_v_0_MPORT_20_data = rf[rf_a_tile_v_0_MPORT_20_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_0_tile_v_3_MPORT_20_en = handshaked & _GEN_1533;
  assign rf_matrix_b_0_tile_v_3_MPORT_20_addr = 8'h70;
  assign rf_matrix_b_0_tile_v_3_MPORT_20_data = rf[rf_matrix_b_0_tile_v_3_MPORT_20_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_0_tile_v_2_MPORT_20_en = handshaked & _GEN_1533;
  assign rf_matrix_b_0_tile_v_2_MPORT_20_addr = 8'h74;
  assign rf_matrix_b_0_tile_v_2_MPORT_20_data = rf[rf_matrix_b_0_tile_v_2_MPORT_20_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_0_tile_v_1_MPORT_20_en = handshaked & _GEN_1533;
  assign rf_matrix_b_0_tile_v_1_MPORT_20_addr = 8'h78;
  assign rf_matrix_b_0_tile_v_1_MPORT_20_data = rf[rf_matrix_b_0_tile_v_1_MPORT_20_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_0_tile_v_0_MPORT_20_en = handshaked & _GEN_1533;
  assign rf_matrix_b_0_tile_v_0_MPORT_20_addr = 8'h7c;
  assign rf_matrix_b_0_tile_v_0_MPORT_20_data = rf[rf_matrix_b_0_tile_v_0_MPORT_20_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_0_tile_v_3_MPORT_20_en = handshaked & _GEN_1533;
  assign rf_matrix_c_0_tile_v_3_MPORT_20_addr = 8'h90;
  assign rf_matrix_c_0_tile_v_3_MPORT_20_data = rf[rf_matrix_c_0_tile_v_3_MPORT_20_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_0_tile_v_2_MPORT_20_en = handshaked & _GEN_1533;
  assign rf_matrix_c_0_tile_v_2_MPORT_20_addr = 8'h91;
  assign rf_matrix_c_0_tile_v_2_MPORT_20_data = rf[rf_matrix_c_0_tile_v_2_MPORT_20_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_0_tile_v_1_MPORT_20_en = handshaked & _GEN_1533;
  assign rf_matrix_c_0_tile_v_1_MPORT_20_addr = 8'h98;
  assign rf_matrix_c_0_tile_v_1_MPORT_20_data = rf[rf_matrix_c_0_tile_v_1_MPORT_20_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_0_tile_v_0_MPORT_20_en = handshaked & _GEN_1533;
  assign rf_matrix_c_0_tile_v_0_MPORT_20_addr = 8'h99;
  assign rf_matrix_c_0_tile_v_0_MPORT_20_data = rf[rf_matrix_c_0_tile_v_0_MPORT_20_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_3_MPORT_7_en = handshaked & _GEN_1545;
  assign rf_a_tile_v_3_MPORT_7_addr = 8'h3;
  assign rf_a_tile_v_3_MPORT_7_data = rf[rf_a_tile_v_3_MPORT_7_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_2_MPORT_7_en = handshaked & _GEN_1545;
  assign rf_a_tile_v_2_MPORT_7_addr = 8'h7;
  assign rf_a_tile_v_2_MPORT_7_data = rf[rf_a_tile_v_2_MPORT_7_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_1_MPORT_21_en = handshaked & _GEN_1545;
  assign rf_a_tile_v_1_MPORT_21_addr = 8'hb;
  assign rf_a_tile_v_1_MPORT_21_data = rf[rf_a_tile_v_1_MPORT_21_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_0_MPORT_21_en = handshaked & _GEN_1545;
  assign rf_a_tile_v_0_MPORT_21_addr = 8'hf;
  assign rf_a_tile_v_0_MPORT_21_data = rf[rf_a_tile_v_0_MPORT_21_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_0_tile_v_3_MPORT_21_en = handshaked & _GEN_1545;
  assign rf_matrix_b_0_tile_v_3_MPORT_21_addr = 8'h70;
  assign rf_matrix_b_0_tile_v_3_MPORT_21_data = rf[rf_matrix_b_0_tile_v_3_MPORT_21_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_0_tile_v_2_MPORT_21_en = handshaked & _GEN_1545;
  assign rf_matrix_b_0_tile_v_2_MPORT_21_addr = 8'h74;
  assign rf_matrix_b_0_tile_v_2_MPORT_21_data = rf[rf_matrix_b_0_tile_v_2_MPORT_21_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_0_tile_v_1_MPORT_21_en = handshaked & _GEN_1545;
  assign rf_matrix_b_0_tile_v_1_MPORT_21_addr = 8'h78;
  assign rf_matrix_b_0_tile_v_1_MPORT_21_data = rf[rf_matrix_b_0_tile_v_1_MPORT_21_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_0_tile_v_0_MPORT_21_en = handshaked & _GEN_1545;
  assign rf_matrix_b_0_tile_v_0_MPORT_21_addr = 8'h7c;
  assign rf_matrix_b_0_tile_v_0_MPORT_21_data = rf[rf_matrix_b_0_tile_v_0_MPORT_21_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_0_tile_v_3_MPORT_21_en = handshaked & _GEN_1545;
  assign rf_matrix_c_0_tile_v_3_MPORT_21_addr = 8'h81;
  assign rf_matrix_c_0_tile_v_3_MPORT_21_data = rf[rf_matrix_c_0_tile_v_3_MPORT_21_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_0_tile_v_2_MPORT_21_en = handshaked & _GEN_1545;
  assign rf_matrix_c_0_tile_v_2_MPORT_21_addr = 8'h85;
  assign rf_matrix_c_0_tile_v_2_MPORT_21_data = rf[rf_matrix_c_0_tile_v_2_MPORT_21_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_0_tile_v_1_MPORT_21_en = handshaked & _GEN_1545;
  assign rf_matrix_c_0_tile_v_1_MPORT_21_addr = 8'h89;
  assign rf_matrix_c_0_tile_v_1_MPORT_21_data = rf[rf_matrix_c_0_tile_v_1_MPORT_21_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_0_tile_v_0_MPORT_21_en = handshaked & _GEN_1545;
  assign rf_matrix_c_0_tile_v_0_MPORT_21_addr = 8'h8d;
  assign rf_matrix_c_0_tile_v_0_MPORT_21_data = rf[rf_matrix_c_0_tile_v_0_MPORT_21_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_1_MPORT_22_en = handshaked & _GEN_1559;
  assign rf_a_tile_v_1_MPORT_22_addr = 8'h3;
  assign rf_a_tile_v_1_MPORT_22_data = rf[rf_a_tile_v_1_MPORT_22_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_0_MPORT_22_en = handshaked & _GEN_1559;
  assign rf_a_tile_v_0_MPORT_22_addr = 8'h7;
  assign rf_a_tile_v_0_MPORT_22_data = rf[rf_a_tile_v_0_MPORT_22_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_0_tile_v_3_MPORT_22_en = handshaked & _GEN_1559;
  assign rf_matrix_b_0_tile_v_3_MPORT_22_addr = 8'h70;
  assign rf_matrix_b_0_tile_v_3_MPORT_22_data = rf[rf_matrix_b_0_tile_v_3_MPORT_22_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_0_tile_v_2_MPORT_22_en = handshaked & _GEN_1559;
  assign rf_matrix_b_0_tile_v_2_MPORT_22_addr = 8'h74;
  assign rf_matrix_b_0_tile_v_2_MPORT_22_data = rf[rf_matrix_b_0_tile_v_2_MPORT_22_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_0_tile_v_1_MPORT_22_en = handshaked & _GEN_1559;
  assign rf_matrix_b_0_tile_v_1_MPORT_22_addr = 8'h78;
  assign rf_matrix_b_0_tile_v_1_MPORT_22_data = rf[rf_matrix_b_0_tile_v_1_MPORT_22_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_0_tile_v_0_MPORT_22_en = handshaked & _GEN_1559;
  assign rf_matrix_b_0_tile_v_0_MPORT_22_addr = 8'h7c;
  assign rf_matrix_b_0_tile_v_0_MPORT_22_data = rf[rf_matrix_b_0_tile_v_0_MPORT_22_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_0_tile_v_3_MPORT_22_en = handshaked & _GEN_1559;
  assign rf_matrix_c_0_tile_v_3_MPORT_22_addr = 8'h82;
  assign rf_matrix_c_0_tile_v_3_MPORT_22_data = rf[rf_matrix_c_0_tile_v_3_MPORT_22_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_0_tile_v_2_MPORT_22_en = handshaked & _GEN_1559;
  assign rf_matrix_c_0_tile_v_2_MPORT_22_addr = 8'h83;
  assign rf_matrix_c_0_tile_v_2_MPORT_22_data = rf[rf_matrix_c_0_tile_v_2_MPORT_22_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_0_tile_v_1_MPORT_22_en = handshaked & _GEN_1559;
  assign rf_matrix_c_0_tile_v_1_MPORT_22_addr = 8'h8a;
  assign rf_matrix_c_0_tile_v_1_MPORT_22_data = rf[rf_matrix_c_0_tile_v_1_MPORT_22_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_0_tile_v_0_MPORT_22_en = handshaked & _GEN_1559;
  assign rf_matrix_c_0_tile_v_0_MPORT_22_addr = 8'h8b;
  assign rf_matrix_c_0_tile_v_0_MPORT_22_data = rf[rf_matrix_c_0_tile_v_0_MPORT_22_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_1_MPORT_23_en = handshaked & _GEN_1571;
  assign rf_a_tile_v_1_MPORT_23_addr = 8'hb;
  assign rf_a_tile_v_1_MPORT_23_data = rf[rf_a_tile_v_1_MPORT_23_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_0_MPORT_23_en = handshaked & _GEN_1571;
  assign rf_a_tile_v_0_MPORT_23_addr = 8'hf;
  assign rf_a_tile_v_0_MPORT_23_data = rf[rf_a_tile_v_0_MPORT_23_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_0_tile_v_3_MPORT_23_en = handshaked & _GEN_1571;
  assign rf_matrix_b_0_tile_v_3_MPORT_23_addr = 8'h70;
  assign rf_matrix_b_0_tile_v_3_MPORT_23_data = rf[rf_matrix_b_0_tile_v_3_MPORT_23_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_0_tile_v_2_MPORT_23_en = handshaked & _GEN_1571;
  assign rf_matrix_b_0_tile_v_2_MPORT_23_addr = 8'h74;
  assign rf_matrix_b_0_tile_v_2_MPORT_23_data = rf[rf_matrix_b_0_tile_v_2_MPORT_23_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_0_tile_v_1_MPORT_23_en = handshaked & _GEN_1571;
  assign rf_matrix_b_0_tile_v_1_MPORT_23_addr = 8'h78;
  assign rf_matrix_b_0_tile_v_1_MPORT_23_data = rf[rf_matrix_b_0_tile_v_1_MPORT_23_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_0_tile_v_0_MPORT_23_en = handshaked & _GEN_1571;
  assign rf_matrix_b_0_tile_v_0_MPORT_23_addr = 8'h7c;
  assign rf_matrix_b_0_tile_v_0_MPORT_23_data = rf[rf_matrix_b_0_tile_v_0_MPORT_23_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_0_tile_v_3_MPORT_23_en = handshaked & _GEN_1571;
  assign rf_matrix_c_0_tile_v_3_MPORT_23_addr = 8'h92;
  assign rf_matrix_c_0_tile_v_3_MPORT_23_data = rf[rf_matrix_c_0_tile_v_3_MPORT_23_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_0_tile_v_2_MPORT_23_en = handshaked & _GEN_1571;
  assign rf_matrix_c_0_tile_v_2_MPORT_23_addr = 8'h93;
  assign rf_matrix_c_0_tile_v_2_MPORT_23_data = rf[rf_matrix_c_0_tile_v_2_MPORT_23_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_0_tile_v_1_MPORT_23_en = handshaked & _GEN_1571;
  assign rf_matrix_c_0_tile_v_1_MPORT_23_addr = 8'h9a;
  assign rf_matrix_c_0_tile_v_1_MPORT_23_data = rf[rf_matrix_c_0_tile_v_1_MPORT_23_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_0_tile_v_0_MPORT_23_en = handshaked & _GEN_1571;
  assign rf_matrix_c_0_tile_v_0_MPORT_23_addr = 8'h9b;
  assign rf_matrix_c_0_tile_v_0_MPORT_23_data = rf[rf_matrix_c_0_tile_v_0_MPORT_23_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_1_MPORT_24_en = handshaked & _GEN_1276;
  assign rf_a_tile_v_1_MPORT_24_addr = 8'h20;
  assign rf_a_tile_v_1_MPORT_24_data = rf[rf_a_tile_v_1_MPORT_24_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_0_MPORT_24_en = handshaked & _GEN_1276;
  assign rf_a_tile_v_0_MPORT_24_addr = 8'h24;
  assign rf_a_tile_v_0_MPORT_24_data = rf[rf_a_tile_v_0_MPORT_24_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_1_tile_v_3_MPORT_en = handshaked & _GEN_1276;
  assign rf_matrix_b_1_tile_v_3_MPORT_addr = 8'h40;
  assign rf_matrix_b_1_tile_v_3_MPORT_data = rf[rf_matrix_b_1_tile_v_3_MPORT_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_1_tile_v_2_MPORT_en = handshaked & _GEN_1276;
  assign rf_matrix_b_1_tile_v_2_MPORT_addr = 8'h44;
  assign rf_matrix_b_1_tile_v_2_MPORT_data = rf[rf_matrix_b_1_tile_v_2_MPORT_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_1_tile_v_1_MPORT_en = handshaked & _GEN_1276;
  assign rf_matrix_b_1_tile_v_1_MPORT_addr = 8'h48;
  assign rf_matrix_b_1_tile_v_1_MPORT_data = rf[rf_matrix_b_1_tile_v_1_MPORT_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_1_tile_v_0_MPORT_en = handshaked & _GEN_1276;
  assign rf_matrix_b_1_tile_v_0_MPORT_addr = 8'h4c;
  assign rf_matrix_b_1_tile_v_0_MPORT_data = rf[rf_matrix_b_1_tile_v_0_MPORT_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_1_tile_v_3_MPORT_en = handshaked & _GEN_1276;
  assign rf_matrix_c_1_tile_v_3_MPORT_addr = 8'hc0;
  assign rf_matrix_c_1_tile_v_3_MPORT_data = rf[rf_matrix_c_1_tile_v_3_MPORT_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_1_tile_v_2_MPORT_en = handshaked & _GEN_1276;
  assign rf_matrix_c_1_tile_v_2_MPORT_addr = 8'hc1;
  assign rf_matrix_c_1_tile_v_2_MPORT_data = rf[rf_matrix_c_1_tile_v_2_MPORT_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_1_tile_v_1_MPORT_en = handshaked & _GEN_1276;
  assign rf_matrix_c_1_tile_v_1_MPORT_addr = 8'hc8;
  assign rf_matrix_c_1_tile_v_1_MPORT_data = rf[rf_matrix_c_1_tile_v_1_MPORT_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_1_tile_v_0_MPORT_en = handshaked & _GEN_1276;
  assign rf_matrix_c_1_tile_v_0_MPORT_addr = 8'hc9;
  assign rf_matrix_c_1_tile_v_0_MPORT_data = rf[rf_matrix_c_1_tile_v_0_MPORT_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_3_MPORT_8_en = handshaked & _GEN_1291;
  assign rf_a_tile_v_3_MPORT_8_addr = 8'h20;
  assign rf_a_tile_v_3_MPORT_8_data = rf[rf_a_tile_v_3_MPORT_8_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_2_MPORT_8_en = handshaked & _GEN_1291;
  assign rf_a_tile_v_2_MPORT_8_addr = 8'h24;
  assign rf_a_tile_v_2_MPORT_8_data = rf[rf_a_tile_v_2_MPORT_8_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_1_MPORT_25_en = handshaked & _GEN_1291;
  assign rf_a_tile_v_1_MPORT_25_addr = 8'h28;
  assign rf_a_tile_v_1_MPORT_25_data = rf[rf_a_tile_v_1_MPORT_25_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_0_MPORT_25_en = handshaked & _GEN_1291;
  assign rf_a_tile_v_0_MPORT_25_addr = 8'h2c;
  assign rf_a_tile_v_0_MPORT_25_data = rf[rf_a_tile_v_0_MPORT_25_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_1_tile_v_3_MPORT_1_en = handshaked & _GEN_1291;
  assign rf_matrix_b_1_tile_v_3_MPORT_1_addr = 8'h40;
  assign rf_matrix_b_1_tile_v_3_MPORT_1_data = rf[rf_matrix_b_1_tile_v_3_MPORT_1_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_1_tile_v_2_MPORT_1_en = handshaked & _GEN_1291;
  assign rf_matrix_b_1_tile_v_2_MPORT_1_addr = 8'h44;
  assign rf_matrix_b_1_tile_v_2_MPORT_1_data = rf[rf_matrix_b_1_tile_v_2_MPORT_1_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_1_tile_v_1_MPORT_1_en = handshaked & _GEN_1291;
  assign rf_matrix_b_1_tile_v_1_MPORT_1_addr = 8'h48;
  assign rf_matrix_b_1_tile_v_1_MPORT_1_data = rf[rf_matrix_b_1_tile_v_1_MPORT_1_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_1_tile_v_0_MPORT_1_en = handshaked & _GEN_1291;
  assign rf_matrix_b_1_tile_v_0_MPORT_1_addr = 8'h4c;
  assign rf_matrix_b_1_tile_v_0_MPORT_1_data = rf[rf_matrix_b_1_tile_v_0_MPORT_1_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_1_tile_v_3_MPORT_1_en = handshaked & _GEN_1291;
  assign rf_matrix_c_1_tile_v_3_MPORT_1_addr = 8'ha0;
  assign rf_matrix_c_1_tile_v_3_MPORT_1_data = rf[rf_matrix_c_1_tile_v_3_MPORT_1_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_1_tile_v_2_MPORT_1_en = handshaked & _GEN_1291;
  assign rf_matrix_c_1_tile_v_2_MPORT_1_addr = 8'ha4;
  assign rf_matrix_c_1_tile_v_2_MPORT_1_data = rf[rf_matrix_c_1_tile_v_2_MPORT_1_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_1_tile_v_1_MPORT_1_en = handshaked & _GEN_1291;
  assign rf_matrix_c_1_tile_v_1_MPORT_1_addr = 8'ha8;
  assign rf_matrix_c_1_tile_v_1_MPORT_1_data = rf[rf_matrix_c_1_tile_v_1_MPORT_1_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_1_tile_v_0_MPORT_1_en = handshaked & _GEN_1291;
  assign rf_matrix_c_1_tile_v_0_MPORT_1_addr = 8'hac;
  assign rf_matrix_c_1_tile_v_0_MPORT_1_data = rf[rf_matrix_c_1_tile_v_0_MPORT_1_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_1_MPORT_26_en = handshaked & _GEN_1305;
  assign rf_a_tile_v_1_MPORT_26_addr = 8'h28;
  assign rf_a_tile_v_1_MPORT_26_data = rf[rf_a_tile_v_1_MPORT_26_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_0_MPORT_26_en = handshaked & _GEN_1305;
  assign rf_a_tile_v_0_MPORT_26_addr = 8'h2c;
  assign rf_a_tile_v_0_MPORT_26_data = rf[rf_a_tile_v_0_MPORT_26_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_1_tile_v_3_MPORT_2_en = handshaked & _GEN_1305;
  assign rf_matrix_b_1_tile_v_3_MPORT_2_addr = 8'h40;
  assign rf_matrix_b_1_tile_v_3_MPORT_2_data = rf[rf_matrix_b_1_tile_v_3_MPORT_2_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_1_tile_v_2_MPORT_2_en = handshaked & _GEN_1305;
  assign rf_matrix_b_1_tile_v_2_MPORT_2_addr = 8'h44;
  assign rf_matrix_b_1_tile_v_2_MPORT_2_data = rf[rf_matrix_b_1_tile_v_2_MPORT_2_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_1_tile_v_1_MPORT_2_en = handshaked & _GEN_1305;
  assign rf_matrix_b_1_tile_v_1_MPORT_2_addr = 8'h48;
  assign rf_matrix_b_1_tile_v_1_MPORT_2_data = rf[rf_matrix_b_1_tile_v_1_MPORT_2_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_1_tile_v_0_MPORT_2_en = handshaked & _GEN_1305;
  assign rf_matrix_b_1_tile_v_0_MPORT_2_addr = 8'h4c;
  assign rf_matrix_b_1_tile_v_0_MPORT_2_data = rf[rf_matrix_b_1_tile_v_0_MPORT_2_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_1_tile_v_3_MPORT_2_en = handshaked & _GEN_1305;
  assign rf_matrix_c_1_tile_v_3_MPORT_2_addr = 8'hd0;
  assign rf_matrix_c_1_tile_v_3_MPORT_2_data = rf[rf_matrix_c_1_tile_v_3_MPORT_2_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_1_tile_v_2_MPORT_2_en = handshaked & _GEN_1305;
  assign rf_matrix_c_1_tile_v_2_MPORT_2_addr = 8'hd1;
  assign rf_matrix_c_1_tile_v_2_MPORT_2_data = rf[rf_matrix_c_1_tile_v_2_MPORT_2_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_1_tile_v_1_MPORT_2_en = handshaked & _GEN_1305;
  assign rf_matrix_c_1_tile_v_1_MPORT_2_addr = 8'hd8;
  assign rf_matrix_c_1_tile_v_1_MPORT_2_data = rf[rf_matrix_c_1_tile_v_1_MPORT_2_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_1_tile_v_0_MPORT_2_en = handshaked & _GEN_1305;
  assign rf_matrix_c_1_tile_v_0_MPORT_2_addr = 8'hd9;
  assign rf_matrix_c_1_tile_v_0_MPORT_2_data = rf[rf_matrix_c_1_tile_v_0_MPORT_2_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_3_MPORT_9_en = handshaked & _GEN_1317;
  assign rf_a_tile_v_3_MPORT_9_addr = 8'h20;
  assign rf_a_tile_v_3_MPORT_9_data = rf[rf_a_tile_v_3_MPORT_9_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_2_MPORT_9_en = handshaked & _GEN_1317;
  assign rf_a_tile_v_2_MPORT_9_addr = 8'h24;
  assign rf_a_tile_v_2_MPORT_9_data = rf[rf_a_tile_v_2_MPORT_9_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_1_MPORT_27_en = handshaked & _GEN_1317;
  assign rf_a_tile_v_1_MPORT_27_addr = 8'h28;
  assign rf_a_tile_v_1_MPORT_27_data = rf[rf_a_tile_v_1_MPORT_27_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_0_MPORT_27_en = handshaked & _GEN_1317;
  assign rf_a_tile_v_0_MPORT_27_addr = 8'h2c;
  assign rf_a_tile_v_0_MPORT_27_data = rf[rf_a_tile_v_0_MPORT_27_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_1_tile_v_3_MPORT_3_en = handshaked & _GEN_1317;
  assign rf_matrix_b_1_tile_v_3_MPORT_3_addr = 8'h40;
  assign rf_matrix_b_1_tile_v_3_MPORT_3_data = rf[rf_matrix_b_1_tile_v_3_MPORT_3_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_1_tile_v_2_MPORT_3_en = handshaked & _GEN_1317;
  assign rf_matrix_b_1_tile_v_2_MPORT_3_addr = 8'h44;
  assign rf_matrix_b_1_tile_v_2_MPORT_3_data = rf[rf_matrix_b_1_tile_v_2_MPORT_3_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_1_tile_v_1_MPORT_3_en = handshaked & _GEN_1317;
  assign rf_matrix_b_1_tile_v_1_MPORT_3_addr = 8'h48;
  assign rf_matrix_b_1_tile_v_1_MPORT_3_data = rf[rf_matrix_b_1_tile_v_1_MPORT_3_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_1_tile_v_0_MPORT_3_en = handshaked & _GEN_1317;
  assign rf_matrix_b_1_tile_v_0_MPORT_3_addr = 8'h4c;
  assign rf_matrix_b_1_tile_v_0_MPORT_3_data = rf[rf_matrix_b_1_tile_v_0_MPORT_3_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_1_tile_v_3_MPORT_3_en = handshaked & _GEN_1317;
  assign rf_matrix_c_1_tile_v_3_MPORT_3_addr = 8'ha1;
  assign rf_matrix_c_1_tile_v_3_MPORT_3_data = rf[rf_matrix_c_1_tile_v_3_MPORT_3_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_1_tile_v_2_MPORT_3_en = handshaked & _GEN_1317;
  assign rf_matrix_c_1_tile_v_2_MPORT_3_addr = 8'ha5;
  assign rf_matrix_c_1_tile_v_2_MPORT_3_data = rf[rf_matrix_c_1_tile_v_2_MPORT_3_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_1_tile_v_1_MPORT_3_en = handshaked & _GEN_1317;
  assign rf_matrix_c_1_tile_v_1_MPORT_3_addr = 8'ha9;
  assign rf_matrix_c_1_tile_v_1_MPORT_3_data = rf[rf_matrix_c_1_tile_v_1_MPORT_3_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_1_tile_v_0_MPORT_3_en = handshaked & _GEN_1317;
  assign rf_matrix_c_1_tile_v_0_MPORT_3_addr = 8'had;
  assign rf_matrix_c_1_tile_v_0_MPORT_3_data = rf[rf_matrix_c_1_tile_v_0_MPORT_3_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_1_MPORT_28_en = handshaked & _GEN_1331;
  assign rf_a_tile_v_1_MPORT_28_addr = 8'h20;
  assign rf_a_tile_v_1_MPORT_28_data = rf[rf_a_tile_v_1_MPORT_28_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_0_MPORT_28_en = handshaked & _GEN_1331;
  assign rf_a_tile_v_0_MPORT_28_addr = 8'h24;
  assign rf_a_tile_v_0_MPORT_28_data = rf[rf_a_tile_v_0_MPORT_28_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_1_tile_v_3_MPORT_4_en = handshaked & _GEN_1331;
  assign rf_matrix_b_1_tile_v_3_MPORT_4_addr = 8'h40;
  assign rf_matrix_b_1_tile_v_3_MPORT_4_data = rf[rf_matrix_b_1_tile_v_3_MPORT_4_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_1_tile_v_2_MPORT_4_en = handshaked & _GEN_1331;
  assign rf_matrix_b_1_tile_v_2_MPORT_4_addr = 8'h44;
  assign rf_matrix_b_1_tile_v_2_MPORT_4_data = rf[rf_matrix_b_1_tile_v_2_MPORT_4_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_1_tile_v_1_MPORT_4_en = handshaked & _GEN_1331;
  assign rf_matrix_b_1_tile_v_1_MPORT_4_addr = 8'h48;
  assign rf_matrix_b_1_tile_v_1_MPORT_4_data = rf[rf_matrix_b_1_tile_v_1_MPORT_4_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_1_tile_v_0_MPORT_4_en = handshaked & _GEN_1331;
  assign rf_matrix_b_1_tile_v_0_MPORT_4_addr = 8'h4c;
  assign rf_matrix_b_1_tile_v_0_MPORT_4_data = rf[rf_matrix_b_1_tile_v_0_MPORT_4_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_1_tile_v_3_MPORT_4_en = handshaked & _GEN_1331;
  assign rf_matrix_c_1_tile_v_3_MPORT_4_addr = 8'hc2;
  assign rf_matrix_c_1_tile_v_3_MPORT_4_data = rf[rf_matrix_c_1_tile_v_3_MPORT_4_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_1_tile_v_2_MPORT_4_en = handshaked & _GEN_1331;
  assign rf_matrix_c_1_tile_v_2_MPORT_4_addr = 8'hc3;
  assign rf_matrix_c_1_tile_v_2_MPORT_4_data = rf[rf_matrix_c_1_tile_v_2_MPORT_4_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_1_tile_v_1_MPORT_4_en = handshaked & _GEN_1331;
  assign rf_matrix_c_1_tile_v_1_MPORT_4_addr = 8'hca;
  assign rf_matrix_c_1_tile_v_1_MPORT_4_data = rf[rf_matrix_c_1_tile_v_1_MPORT_4_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_1_tile_v_0_MPORT_4_en = handshaked & _GEN_1331;
  assign rf_matrix_c_1_tile_v_0_MPORT_4_addr = 8'hcb;
  assign rf_matrix_c_1_tile_v_0_MPORT_4_data = rf[rf_matrix_c_1_tile_v_0_MPORT_4_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_1_MPORT_29_en = handshaked & _GEN_1343;
  assign rf_a_tile_v_1_MPORT_29_addr = 8'h28;
  assign rf_a_tile_v_1_MPORT_29_data = rf[rf_a_tile_v_1_MPORT_29_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_0_MPORT_29_en = handshaked & _GEN_1343;
  assign rf_a_tile_v_0_MPORT_29_addr = 8'h2c;
  assign rf_a_tile_v_0_MPORT_29_data = rf[rf_a_tile_v_0_MPORT_29_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_1_tile_v_3_MPORT_5_en = handshaked & _GEN_1343;
  assign rf_matrix_b_1_tile_v_3_MPORT_5_addr = 8'h40;
  assign rf_matrix_b_1_tile_v_3_MPORT_5_data = rf[rf_matrix_b_1_tile_v_3_MPORT_5_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_1_tile_v_2_MPORT_5_en = handshaked & _GEN_1343;
  assign rf_matrix_b_1_tile_v_2_MPORT_5_addr = 8'h44;
  assign rf_matrix_b_1_tile_v_2_MPORT_5_data = rf[rf_matrix_b_1_tile_v_2_MPORT_5_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_1_tile_v_1_MPORT_5_en = handshaked & _GEN_1343;
  assign rf_matrix_b_1_tile_v_1_MPORT_5_addr = 8'h48;
  assign rf_matrix_b_1_tile_v_1_MPORT_5_data = rf[rf_matrix_b_1_tile_v_1_MPORT_5_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_1_tile_v_0_MPORT_5_en = handshaked & _GEN_1343;
  assign rf_matrix_b_1_tile_v_0_MPORT_5_addr = 8'h4c;
  assign rf_matrix_b_1_tile_v_0_MPORT_5_data = rf[rf_matrix_b_1_tile_v_0_MPORT_5_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_1_tile_v_3_MPORT_5_en = handshaked & _GEN_1343;
  assign rf_matrix_c_1_tile_v_3_MPORT_5_addr = 8'hd2;
  assign rf_matrix_c_1_tile_v_3_MPORT_5_data = rf[rf_matrix_c_1_tile_v_3_MPORT_5_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_1_tile_v_2_MPORT_5_en = handshaked & _GEN_1343;
  assign rf_matrix_c_1_tile_v_2_MPORT_5_addr = 8'hd3;
  assign rf_matrix_c_1_tile_v_2_MPORT_5_data = rf[rf_matrix_c_1_tile_v_2_MPORT_5_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_1_tile_v_1_MPORT_5_en = handshaked & _GEN_1343;
  assign rf_matrix_c_1_tile_v_1_MPORT_5_addr = 8'hda;
  assign rf_matrix_c_1_tile_v_1_MPORT_5_data = rf[rf_matrix_c_1_tile_v_1_MPORT_5_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_1_tile_v_0_MPORT_5_en = handshaked & _GEN_1343;
  assign rf_matrix_c_1_tile_v_0_MPORT_5_addr = 8'hdb;
  assign rf_matrix_c_1_tile_v_0_MPORT_5_data = rf[rf_matrix_c_1_tile_v_0_MPORT_5_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_1_MPORT_30_en = handshaked & _GEN_1355;
  assign rf_a_tile_v_1_MPORT_30_addr = 8'h21;
  assign rf_a_tile_v_1_MPORT_30_data = rf[rf_a_tile_v_1_MPORT_30_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_0_MPORT_30_en = handshaked & _GEN_1355;
  assign rf_a_tile_v_0_MPORT_30_addr = 8'h25;
  assign rf_a_tile_v_0_MPORT_30_data = rf[rf_a_tile_v_0_MPORT_30_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_1_tile_v_3_MPORT_6_en = handshaked & _GEN_1355;
  assign rf_matrix_b_1_tile_v_3_MPORT_6_addr = 8'h50;
  assign rf_matrix_b_1_tile_v_3_MPORT_6_data = rf[rf_matrix_b_1_tile_v_3_MPORT_6_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_1_tile_v_2_MPORT_6_en = handshaked & _GEN_1355;
  assign rf_matrix_b_1_tile_v_2_MPORT_6_addr = 8'h54;
  assign rf_matrix_b_1_tile_v_2_MPORT_6_data = rf[rf_matrix_b_1_tile_v_2_MPORT_6_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_1_tile_v_1_MPORT_6_en = handshaked & _GEN_1355;
  assign rf_matrix_b_1_tile_v_1_MPORT_6_addr = 8'h58;
  assign rf_matrix_b_1_tile_v_1_MPORT_6_data = rf[rf_matrix_b_1_tile_v_1_MPORT_6_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_1_tile_v_0_MPORT_6_en = handshaked & _GEN_1355;
  assign rf_matrix_b_1_tile_v_0_MPORT_6_addr = 8'h5c;
  assign rf_matrix_b_1_tile_v_0_MPORT_6_data = rf[rf_matrix_b_1_tile_v_0_MPORT_6_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_1_tile_v_3_MPORT_6_en = handshaked & _GEN_1355;
  assign rf_matrix_c_1_tile_v_3_MPORT_6_addr = 8'hc0;
  assign rf_matrix_c_1_tile_v_3_MPORT_6_data = rf[rf_matrix_c_1_tile_v_3_MPORT_6_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_1_tile_v_2_MPORT_6_en = handshaked & _GEN_1355;
  assign rf_matrix_c_1_tile_v_2_MPORT_6_addr = 8'hc1;
  assign rf_matrix_c_1_tile_v_2_MPORT_6_data = rf[rf_matrix_c_1_tile_v_2_MPORT_6_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_1_tile_v_1_MPORT_6_en = handshaked & _GEN_1355;
  assign rf_matrix_c_1_tile_v_1_MPORT_6_addr = 8'hc8;
  assign rf_matrix_c_1_tile_v_1_MPORT_6_data = rf[rf_matrix_c_1_tile_v_1_MPORT_6_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_1_tile_v_0_MPORT_6_en = handshaked & _GEN_1355;
  assign rf_matrix_c_1_tile_v_0_MPORT_6_addr = 8'hc9;
  assign rf_matrix_c_1_tile_v_0_MPORT_6_data = rf[rf_matrix_c_1_tile_v_0_MPORT_6_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_3_MPORT_10_en = handshaked & _GEN_1367;
  assign rf_a_tile_v_3_MPORT_10_addr = 8'h21;
  assign rf_a_tile_v_3_MPORT_10_data = rf[rf_a_tile_v_3_MPORT_10_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_2_MPORT_10_en = handshaked & _GEN_1367;
  assign rf_a_tile_v_2_MPORT_10_addr = 8'h25;
  assign rf_a_tile_v_2_MPORT_10_data = rf[rf_a_tile_v_2_MPORT_10_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_1_MPORT_31_en = handshaked & _GEN_1367;
  assign rf_a_tile_v_1_MPORT_31_addr = 8'h29;
  assign rf_a_tile_v_1_MPORT_31_data = rf[rf_a_tile_v_1_MPORT_31_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_0_MPORT_31_en = handshaked & _GEN_1367;
  assign rf_a_tile_v_0_MPORT_31_addr = 8'h2d;
  assign rf_a_tile_v_0_MPORT_31_data = rf[rf_a_tile_v_0_MPORT_31_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_1_tile_v_3_MPORT_7_en = handshaked & _GEN_1367;
  assign rf_matrix_b_1_tile_v_3_MPORT_7_addr = 8'h50;
  assign rf_matrix_b_1_tile_v_3_MPORT_7_data = rf[rf_matrix_b_1_tile_v_3_MPORT_7_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_1_tile_v_2_MPORT_7_en = handshaked & _GEN_1367;
  assign rf_matrix_b_1_tile_v_2_MPORT_7_addr = 8'h54;
  assign rf_matrix_b_1_tile_v_2_MPORT_7_data = rf[rf_matrix_b_1_tile_v_2_MPORT_7_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_1_tile_v_1_MPORT_7_en = handshaked & _GEN_1367;
  assign rf_matrix_b_1_tile_v_1_MPORT_7_addr = 8'h58;
  assign rf_matrix_b_1_tile_v_1_MPORT_7_data = rf[rf_matrix_b_1_tile_v_1_MPORT_7_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_1_tile_v_0_MPORT_7_en = handshaked & _GEN_1367;
  assign rf_matrix_b_1_tile_v_0_MPORT_7_addr = 8'h5c;
  assign rf_matrix_b_1_tile_v_0_MPORT_7_data = rf[rf_matrix_b_1_tile_v_0_MPORT_7_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_1_tile_v_3_MPORT_7_en = handshaked & _GEN_1367;
  assign rf_matrix_c_1_tile_v_3_MPORT_7_addr = 8'ha0;
  assign rf_matrix_c_1_tile_v_3_MPORT_7_data = rf[rf_matrix_c_1_tile_v_3_MPORT_7_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_1_tile_v_2_MPORT_7_en = handshaked & _GEN_1367;
  assign rf_matrix_c_1_tile_v_2_MPORT_7_addr = 8'ha4;
  assign rf_matrix_c_1_tile_v_2_MPORT_7_data = rf[rf_matrix_c_1_tile_v_2_MPORT_7_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_1_tile_v_1_MPORT_7_en = handshaked & _GEN_1367;
  assign rf_matrix_c_1_tile_v_1_MPORT_7_addr = 8'ha8;
  assign rf_matrix_c_1_tile_v_1_MPORT_7_data = rf[rf_matrix_c_1_tile_v_1_MPORT_7_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_1_tile_v_0_MPORT_7_en = handshaked & _GEN_1367;
  assign rf_matrix_c_1_tile_v_0_MPORT_7_addr = 8'hac;
  assign rf_matrix_c_1_tile_v_0_MPORT_7_data = rf[rf_matrix_c_1_tile_v_0_MPORT_7_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_1_MPORT_32_en = handshaked & _GEN_1381;
  assign rf_a_tile_v_1_MPORT_32_addr = 8'h29;
  assign rf_a_tile_v_1_MPORT_32_data = rf[rf_a_tile_v_1_MPORT_32_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_0_MPORT_32_en = handshaked & _GEN_1381;
  assign rf_a_tile_v_0_MPORT_32_addr = 8'h2d;
  assign rf_a_tile_v_0_MPORT_32_data = rf[rf_a_tile_v_0_MPORT_32_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_1_tile_v_3_MPORT_8_en = handshaked & _GEN_1381;
  assign rf_matrix_b_1_tile_v_3_MPORT_8_addr = 8'h50;
  assign rf_matrix_b_1_tile_v_3_MPORT_8_data = rf[rf_matrix_b_1_tile_v_3_MPORT_8_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_1_tile_v_2_MPORT_8_en = handshaked & _GEN_1381;
  assign rf_matrix_b_1_tile_v_2_MPORT_8_addr = 8'h54;
  assign rf_matrix_b_1_tile_v_2_MPORT_8_data = rf[rf_matrix_b_1_tile_v_2_MPORT_8_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_1_tile_v_1_MPORT_8_en = handshaked & _GEN_1381;
  assign rf_matrix_b_1_tile_v_1_MPORT_8_addr = 8'h58;
  assign rf_matrix_b_1_tile_v_1_MPORT_8_data = rf[rf_matrix_b_1_tile_v_1_MPORT_8_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_1_tile_v_0_MPORT_8_en = handshaked & _GEN_1381;
  assign rf_matrix_b_1_tile_v_0_MPORT_8_addr = 8'h5c;
  assign rf_matrix_b_1_tile_v_0_MPORT_8_data = rf[rf_matrix_b_1_tile_v_0_MPORT_8_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_1_tile_v_3_MPORT_8_en = handshaked & _GEN_1381;
  assign rf_matrix_c_1_tile_v_3_MPORT_8_addr = 8'hd0;
  assign rf_matrix_c_1_tile_v_3_MPORT_8_data = rf[rf_matrix_c_1_tile_v_3_MPORT_8_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_1_tile_v_2_MPORT_8_en = handshaked & _GEN_1381;
  assign rf_matrix_c_1_tile_v_2_MPORT_8_addr = 8'hd1;
  assign rf_matrix_c_1_tile_v_2_MPORT_8_data = rf[rf_matrix_c_1_tile_v_2_MPORT_8_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_1_tile_v_1_MPORT_8_en = handshaked & _GEN_1381;
  assign rf_matrix_c_1_tile_v_1_MPORT_8_addr = 8'hd8;
  assign rf_matrix_c_1_tile_v_1_MPORT_8_data = rf[rf_matrix_c_1_tile_v_1_MPORT_8_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_1_tile_v_0_MPORT_8_en = handshaked & _GEN_1381;
  assign rf_matrix_c_1_tile_v_0_MPORT_8_addr = 8'hd9;
  assign rf_matrix_c_1_tile_v_0_MPORT_8_data = rf[rf_matrix_c_1_tile_v_0_MPORT_8_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_3_MPORT_11_en = handshaked & _GEN_1393;
  assign rf_a_tile_v_3_MPORT_11_addr = 8'h21;
  assign rf_a_tile_v_3_MPORT_11_data = rf[rf_a_tile_v_3_MPORT_11_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_2_MPORT_11_en = handshaked & _GEN_1393;
  assign rf_a_tile_v_2_MPORT_11_addr = 8'h25;
  assign rf_a_tile_v_2_MPORT_11_data = rf[rf_a_tile_v_2_MPORT_11_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_1_MPORT_33_en = handshaked & _GEN_1393;
  assign rf_a_tile_v_1_MPORT_33_addr = 8'h29;
  assign rf_a_tile_v_1_MPORT_33_data = rf[rf_a_tile_v_1_MPORT_33_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_0_MPORT_33_en = handshaked & _GEN_1393;
  assign rf_a_tile_v_0_MPORT_33_addr = 8'h2d;
  assign rf_a_tile_v_0_MPORT_33_data = rf[rf_a_tile_v_0_MPORT_33_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_1_tile_v_3_MPORT_9_en = handshaked & _GEN_1393;
  assign rf_matrix_b_1_tile_v_3_MPORT_9_addr = 8'h50;
  assign rf_matrix_b_1_tile_v_3_MPORT_9_data = rf[rf_matrix_b_1_tile_v_3_MPORT_9_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_1_tile_v_2_MPORT_9_en = handshaked & _GEN_1393;
  assign rf_matrix_b_1_tile_v_2_MPORT_9_addr = 8'h54;
  assign rf_matrix_b_1_tile_v_2_MPORT_9_data = rf[rf_matrix_b_1_tile_v_2_MPORT_9_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_1_tile_v_1_MPORT_9_en = handshaked & _GEN_1393;
  assign rf_matrix_b_1_tile_v_1_MPORT_9_addr = 8'h58;
  assign rf_matrix_b_1_tile_v_1_MPORT_9_data = rf[rf_matrix_b_1_tile_v_1_MPORT_9_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_1_tile_v_0_MPORT_9_en = handshaked & _GEN_1393;
  assign rf_matrix_b_1_tile_v_0_MPORT_9_addr = 8'h5c;
  assign rf_matrix_b_1_tile_v_0_MPORT_9_data = rf[rf_matrix_b_1_tile_v_0_MPORT_9_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_1_tile_v_3_MPORT_9_en = handshaked & _GEN_1393;
  assign rf_matrix_c_1_tile_v_3_MPORT_9_addr = 8'ha1;
  assign rf_matrix_c_1_tile_v_3_MPORT_9_data = rf[rf_matrix_c_1_tile_v_3_MPORT_9_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_1_tile_v_2_MPORT_9_en = handshaked & _GEN_1393;
  assign rf_matrix_c_1_tile_v_2_MPORT_9_addr = 8'ha5;
  assign rf_matrix_c_1_tile_v_2_MPORT_9_data = rf[rf_matrix_c_1_tile_v_2_MPORT_9_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_1_tile_v_1_MPORT_9_en = handshaked & _GEN_1393;
  assign rf_matrix_c_1_tile_v_1_MPORT_9_addr = 8'ha9;
  assign rf_matrix_c_1_tile_v_1_MPORT_9_data = rf[rf_matrix_c_1_tile_v_1_MPORT_9_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_1_tile_v_0_MPORT_9_en = handshaked & _GEN_1393;
  assign rf_matrix_c_1_tile_v_0_MPORT_9_addr = 8'had;
  assign rf_matrix_c_1_tile_v_0_MPORT_9_data = rf[rf_matrix_c_1_tile_v_0_MPORT_9_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_1_MPORT_34_en = handshaked & _GEN_1407;
  assign rf_a_tile_v_1_MPORT_34_addr = 8'h21;
  assign rf_a_tile_v_1_MPORT_34_data = rf[rf_a_tile_v_1_MPORT_34_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_0_MPORT_34_en = handshaked & _GEN_1407;
  assign rf_a_tile_v_0_MPORT_34_addr = 8'h25;
  assign rf_a_tile_v_0_MPORT_34_data = rf[rf_a_tile_v_0_MPORT_34_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_1_tile_v_3_MPORT_10_en = handshaked & _GEN_1407;
  assign rf_matrix_b_1_tile_v_3_MPORT_10_addr = 8'h50;
  assign rf_matrix_b_1_tile_v_3_MPORT_10_data = rf[rf_matrix_b_1_tile_v_3_MPORT_10_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_1_tile_v_2_MPORT_10_en = handshaked & _GEN_1407;
  assign rf_matrix_b_1_tile_v_2_MPORT_10_addr = 8'h54;
  assign rf_matrix_b_1_tile_v_2_MPORT_10_data = rf[rf_matrix_b_1_tile_v_2_MPORT_10_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_1_tile_v_1_MPORT_10_en = handshaked & _GEN_1407;
  assign rf_matrix_b_1_tile_v_1_MPORT_10_addr = 8'h58;
  assign rf_matrix_b_1_tile_v_1_MPORT_10_data = rf[rf_matrix_b_1_tile_v_1_MPORT_10_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_1_tile_v_0_MPORT_10_en = handshaked & _GEN_1407;
  assign rf_matrix_b_1_tile_v_0_MPORT_10_addr = 8'h5c;
  assign rf_matrix_b_1_tile_v_0_MPORT_10_data = rf[rf_matrix_b_1_tile_v_0_MPORT_10_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_1_tile_v_3_MPORT_10_en = handshaked & _GEN_1407;
  assign rf_matrix_c_1_tile_v_3_MPORT_10_addr = 8'hc2;
  assign rf_matrix_c_1_tile_v_3_MPORT_10_data = rf[rf_matrix_c_1_tile_v_3_MPORT_10_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_1_tile_v_2_MPORT_10_en = handshaked & _GEN_1407;
  assign rf_matrix_c_1_tile_v_2_MPORT_10_addr = 8'hc3;
  assign rf_matrix_c_1_tile_v_2_MPORT_10_data = rf[rf_matrix_c_1_tile_v_2_MPORT_10_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_1_tile_v_1_MPORT_10_en = handshaked & _GEN_1407;
  assign rf_matrix_c_1_tile_v_1_MPORT_10_addr = 8'hca;
  assign rf_matrix_c_1_tile_v_1_MPORT_10_data = rf[rf_matrix_c_1_tile_v_1_MPORT_10_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_1_tile_v_0_MPORT_10_en = handshaked & _GEN_1407;
  assign rf_matrix_c_1_tile_v_0_MPORT_10_addr = 8'hcb;
  assign rf_matrix_c_1_tile_v_0_MPORT_10_data = rf[rf_matrix_c_1_tile_v_0_MPORT_10_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_1_MPORT_35_en = handshaked & _GEN_1419;
  assign rf_a_tile_v_1_MPORT_35_addr = 8'h29;
  assign rf_a_tile_v_1_MPORT_35_data = rf[rf_a_tile_v_1_MPORT_35_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_0_MPORT_35_en = handshaked & _GEN_1419;
  assign rf_a_tile_v_0_MPORT_35_addr = 8'h2d;
  assign rf_a_tile_v_0_MPORT_35_data = rf[rf_a_tile_v_0_MPORT_35_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_1_tile_v_3_MPORT_11_en = handshaked & _GEN_1419;
  assign rf_matrix_b_1_tile_v_3_MPORT_11_addr = 8'h50;
  assign rf_matrix_b_1_tile_v_3_MPORT_11_data = rf[rf_matrix_b_1_tile_v_3_MPORT_11_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_1_tile_v_2_MPORT_11_en = handshaked & _GEN_1419;
  assign rf_matrix_b_1_tile_v_2_MPORT_11_addr = 8'h54;
  assign rf_matrix_b_1_tile_v_2_MPORT_11_data = rf[rf_matrix_b_1_tile_v_2_MPORT_11_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_1_tile_v_1_MPORT_11_en = handshaked & _GEN_1419;
  assign rf_matrix_b_1_tile_v_1_MPORT_11_addr = 8'h58;
  assign rf_matrix_b_1_tile_v_1_MPORT_11_data = rf[rf_matrix_b_1_tile_v_1_MPORT_11_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_1_tile_v_0_MPORT_11_en = handshaked & _GEN_1419;
  assign rf_matrix_b_1_tile_v_0_MPORT_11_addr = 8'h5c;
  assign rf_matrix_b_1_tile_v_0_MPORT_11_data = rf[rf_matrix_b_1_tile_v_0_MPORT_11_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_1_tile_v_3_MPORT_11_en = handshaked & _GEN_1419;
  assign rf_matrix_c_1_tile_v_3_MPORT_11_addr = 8'hd2;
  assign rf_matrix_c_1_tile_v_3_MPORT_11_data = rf[rf_matrix_c_1_tile_v_3_MPORT_11_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_1_tile_v_2_MPORT_11_en = handshaked & _GEN_1419;
  assign rf_matrix_c_1_tile_v_2_MPORT_11_addr = 8'hd3;
  assign rf_matrix_c_1_tile_v_2_MPORT_11_data = rf[rf_matrix_c_1_tile_v_2_MPORT_11_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_1_tile_v_1_MPORT_11_en = handshaked & _GEN_1419;
  assign rf_matrix_c_1_tile_v_1_MPORT_11_addr = 8'hda;
  assign rf_matrix_c_1_tile_v_1_MPORT_11_data = rf[rf_matrix_c_1_tile_v_1_MPORT_11_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_1_tile_v_0_MPORT_11_en = handshaked & _GEN_1419;
  assign rf_matrix_c_1_tile_v_0_MPORT_11_addr = 8'hdb;
  assign rf_matrix_c_1_tile_v_0_MPORT_11_data = rf[rf_matrix_c_1_tile_v_0_MPORT_11_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_1_MPORT_36_en = handshaked & _GEN_1431;
  assign rf_a_tile_v_1_MPORT_36_addr = 8'h22;
  assign rf_a_tile_v_1_MPORT_36_data = rf[rf_a_tile_v_1_MPORT_36_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_0_MPORT_36_en = handshaked & _GEN_1431;
  assign rf_a_tile_v_0_MPORT_36_addr = 8'h26;
  assign rf_a_tile_v_0_MPORT_36_data = rf[rf_a_tile_v_0_MPORT_36_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_1_tile_v_3_MPORT_12_en = handshaked & _GEN_1431;
  assign rf_matrix_b_1_tile_v_3_MPORT_12_addr = 8'h60;
  assign rf_matrix_b_1_tile_v_3_MPORT_12_data = rf[rf_matrix_b_1_tile_v_3_MPORT_12_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_1_tile_v_2_MPORT_12_en = handshaked & _GEN_1431;
  assign rf_matrix_b_1_tile_v_2_MPORT_12_addr = 8'h64;
  assign rf_matrix_b_1_tile_v_2_MPORT_12_data = rf[rf_matrix_b_1_tile_v_2_MPORT_12_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_1_tile_v_1_MPORT_12_en = handshaked & _GEN_1431;
  assign rf_matrix_b_1_tile_v_1_MPORT_12_addr = 8'h68;
  assign rf_matrix_b_1_tile_v_1_MPORT_12_data = rf[rf_matrix_b_1_tile_v_1_MPORT_12_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_1_tile_v_0_MPORT_12_en = handshaked & _GEN_1431;
  assign rf_matrix_b_1_tile_v_0_MPORT_12_addr = 8'h6c;
  assign rf_matrix_b_1_tile_v_0_MPORT_12_data = rf[rf_matrix_b_1_tile_v_0_MPORT_12_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_1_tile_v_3_MPORT_12_en = handshaked & _GEN_1431;
  assign rf_matrix_c_1_tile_v_3_MPORT_12_addr = 8'hc0;
  assign rf_matrix_c_1_tile_v_3_MPORT_12_data = rf[rf_matrix_c_1_tile_v_3_MPORT_12_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_1_tile_v_2_MPORT_12_en = handshaked & _GEN_1431;
  assign rf_matrix_c_1_tile_v_2_MPORT_12_addr = 8'hc1;
  assign rf_matrix_c_1_tile_v_2_MPORT_12_data = rf[rf_matrix_c_1_tile_v_2_MPORT_12_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_1_tile_v_1_MPORT_12_en = handshaked & _GEN_1431;
  assign rf_matrix_c_1_tile_v_1_MPORT_12_addr = 8'hc8;
  assign rf_matrix_c_1_tile_v_1_MPORT_12_data = rf[rf_matrix_c_1_tile_v_1_MPORT_12_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_1_tile_v_0_MPORT_12_en = handshaked & _GEN_1431;
  assign rf_matrix_c_1_tile_v_0_MPORT_12_addr = 8'hc9;
  assign rf_matrix_c_1_tile_v_0_MPORT_12_data = rf[rf_matrix_c_1_tile_v_0_MPORT_12_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_3_MPORT_12_en = handshaked & _GEN_1443;
  assign rf_a_tile_v_3_MPORT_12_addr = 8'h22;
  assign rf_a_tile_v_3_MPORT_12_data = rf[rf_a_tile_v_3_MPORT_12_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_2_MPORT_12_en = handshaked & _GEN_1443;
  assign rf_a_tile_v_2_MPORT_12_addr = 8'h26;
  assign rf_a_tile_v_2_MPORT_12_data = rf[rf_a_tile_v_2_MPORT_12_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_1_MPORT_37_en = handshaked & _GEN_1443;
  assign rf_a_tile_v_1_MPORT_37_addr = 8'h2a;
  assign rf_a_tile_v_1_MPORT_37_data = rf[rf_a_tile_v_1_MPORT_37_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_0_MPORT_37_en = handshaked & _GEN_1443;
  assign rf_a_tile_v_0_MPORT_37_addr = 8'h2e;
  assign rf_a_tile_v_0_MPORT_37_data = rf[rf_a_tile_v_0_MPORT_37_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_1_tile_v_3_MPORT_13_en = handshaked & _GEN_1443;
  assign rf_matrix_b_1_tile_v_3_MPORT_13_addr = 8'h60;
  assign rf_matrix_b_1_tile_v_3_MPORT_13_data = rf[rf_matrix_b_1_tile_v_3_MPORT_13_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_1_tile_v_2_MPORT_13_en = handshaked & _GEN_1443;
  assign rf_matrix_b_1_tile_v_2_MPORT_13_addr = 8'h64;
  assign rf_matrix_b_1_tile_v_2_MPORT_13_data = rf[rf_matrix_b_1_tile_v_2_MPORT_13_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_1_tile_v_1_MPORT_13_en = handshaked & _GEN_1443;
  assign rf_matrix_b_1_tile_v_1_MPORT_13_addr = 8'h68;
  assign rf_matrix_b_1_tile_v_1_MPORT_13_data = rf[rf_matrix_b_1_tile_v_1_MPORT_13_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_1_tile_v_0_MPORT_13_en = handshaked & _GEN_1443;
  assign rf_matrix_b_1_tile_v_0_MPORT_13_addr = 8'h6c;
  assign rf_matrix_b_1_tile_v_0_MPORT_13_data = rf[rf_matrix_b_1_tile_v_0_MPORT_13_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_1_tile_v_3_MPORT_13_en = handshaked & _GEN_1443;
  assign rf_matrix_c_1_tile_v_3_MPORT_13_addr = 8'ha0;
  assign rf_matrix_c_1_tile_v_3_MPORT_13_data = rf[rf_matrix_c_1_tile_v_3_MPORT_13_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_1_tile_v_2_MPORT_13_en = handshaked & _GEN_1443;
  assign rf_matrix_c_1_tile_v_2_MPORT_13_addr = 8'ha4;
  assign rf_matrix_c_1_tile_v_2_MPORT_13_data = rf[rf_matrix_c_1_tile_v_2_MPORT_13_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_1_tile_v_1_MPORT_13_en = handshaked & _GEN_1443;
  assign rf_matrix_c_1_tile_v_1_MPORT_13_addr = 8'ha8;
  assign rf_matrix_c_1_tile_v_1_MPORT_13_data = rf[rf_matrix_c_1_tile_v_1_MPORT_13_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_1_tile_v_0_MPORT_13_en = handshaked & _GEN_1443;
  assign rf_matrix_c_1_tile_v_0_MPORT_13_addr = 8'hac;
  assign rf_matrix_c_1_tile_v_0_MPORT_13_data = rf[rf_matrix_c_1_tile_v_0_MPORT_13_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_1_MPORT_38_en = handshaked & _GEN_1457;
  assign rf_a_tile_v_1_MPORT_38_addr = 8'h2a;
  assign rf_a_tile_v_1_MPORT_38_data = rf[rf_a_tile_v_1_MPORT_38_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_0_MPORT_38_en = handshaked & _GEN_1457;
  assign rf_a_tile_v_0_MPORT_38_addr = 8'h2e;
  assign rf_a_tile_v_0_MPORT_38_data = rf[rf_a_tile_v_0_MPORT_38_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_1_tile_v_3_MPORT_14_en = handshaked & _GEN_1457;
  assign rf_matrix_b_1_tile_v_3_MPORT_14_addr = 8'h60;
  assign rf_matrix_b_1_tile_v_3_MPORT_14_data = rf[rf_matrix_b_1_tile_v_3_MPORT_14_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_1_tile_v_2_MPORT_14_en = handshaked & _GEN_1457;
  assign rf_matrix_b_1_tile_v_2_MPORT_14_addr = 8'h64;
  assign rf_matrix_b_1_tile_v_2_MPORT_14_data = rf[rf_matrix_b_1_tile_v_2_MPORT_14_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_1_tile_v_1_MPORT_14_en = handshaked & _GEN_1457;
  assign rf_matrix_b_1_tile_v_1_MPORT_14_addr = 8'h68;
  assign rf_matrix_b_1_tile_v_1_MPORT_14_data = rf[rf_matrix_b_1_tile_v_1_MPORT_14_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_1_tile_v_0_MPORT_14_en = handshaked & _GEN_1457;
  assign rf_matrix_b_1_tile_v_0_MPORT_14_addr = 8'h6c;
  assign rf_matrix_b_1_tile_v_0_MPORT_14_data = rf[rf_matrix_b_1_tile_v_0_MPORT_14_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_1_tile_v_3_MPORT_14_en = handshaked & _GEN_1457;
  assign rf_matrix_c_1_tile_v_3_MPORT_14_addr = 8'hd0;
  assign rf_matrix_c_1_tile_v_3_MPORT_14_data = rf[rf_matrix_c_1_tile_v_3_MPORT_14_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_1_tile_v_2_MPORT_14_en = handshaked & _GEN_1457;
  assign rf_matrix_c_1_tile_v_2_MPORT_14_addr = 8'hd1;
  assign rf_matrix_c_1_tile_v_2_MPORT_14_data = rf[rf_matrix_c_1_tile_v_2_MPORT_14_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_1_tile_v_1_MPORT_14_en = handshaked & _GEN_1457;
  assign rf_matrix_c_1_tile_v_1_MPORT_14_addr = 8'hd8;
  assign rf_matrix_c_1_tile_v_1_MPORT_14_data = rf[rf_matrix_c_1_tile_v_1_MPORT_14_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_1_tile_v_0_MPORT_14_en = handshaked & _GEN_1457;
  assign rf_matrix_c_1_tile_v_0_MPORT_14_addr = 8'hd9;
  assign rf_matrix_c_1_tile_v_0_MPORT_14_data = rf[rf_matrix_c_1_tile_v_0_MPORT_14_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_3_MPORT_13_en = handshaked & _GEN_1469;
  assign rf_a_tile_v_3_MPORT_13_addr = 8'h22;
  assign rf_a_tile_v_3_MPORT_13_data = rf[rf_a_tile_v_3_MPORT_13_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_2_MPORT_13_en = handshaked & _GEN_1469;
  assign rf_a_tile_v_2_MPORT_13_addr = 8'h26;
  assign rf_a_tile_v_2_MPORT_13_data = rf[rf_a_tile_v_2_MPORT_13_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_1_MPORT_39_en = handshaked & _GEN_1469;
  assign rf_a_tile_v_1_MPORT_39_addr = 8'h2a;
  assign rf_a_tile_v_1_MPORT_39_data = rf[rf_a_tile_v_1_MPORT_39_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_0_MPORT_39_en = handshaked & _GEN_1469;
  assign rf_a_tile_v_0_MPORT_39_addr = 8'h2e;
  assign rf_a_tile_v_0_MPORT_39_data = rf[rf_a_tile_v_0_MPORT_39_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_1_tile_v_3_MPORT_15_en = handshaked & _GEN_1469;
  assign rf_matrix_b_1_tile_v_3_MPORT_15_addr = 8'h60;
  assign rf_matrix_b_1_tile_v_3_MPORT_15_data = rf[rf_matrix_b_1_tile_v_3_MPORT_15_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_1_tile_v_2_MPORT_15_en = handshaked & _GEN_1469;
  assign rf_matrix_b_1_tile_v_2_MPORT_15_addr = 8'h64;
  assign rf_matrix_b_1_tile_v_2_MPORT_15_data = rf[rf_matrix_b_1_tile_v_2_MPORT_15_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_1_tile_v_1_MPORT_15_en = handshaked & _GEN_1469;
  assign rf_matrix_b_1_tile_v_1_MPORT_15_addr = 8'h68;
  assign rf_matrix_b_1_tile_v_1_MPORT_15_data = rf[rf_matrix_b_1_tile_v_1_MPORT_15_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_1_tile_v_0_MPORT_15_en = handshaked & _GEN_1469;
  assign rf_matrix_b_1_tile_v_0_MPORT_15_addr = 8'h6c;
  assign rf_matrix_b_1_tile_v_0_MPORT_15_data = rf[rf_matrix_b_1_tile_v_0_MPORT_15_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_1_tile_v_3_MPORT_15_en = handshaked & _GEN_1469;
  assign rf_matrix_c_1_tile_v_3_MPORT_15_addr = 8'ha1;
  assign rf_matrix_c_1_tile_v_3_MPORT_15_data = rf[rf_matrix_c_1_tile_v_3_MPORT_15_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_1_tile_v_2_MPORT_15_en = handshaked & _GEN_1469;
  assign rf_matrix_c_1_tile_v_2_MPORT_15_addr = 8'ha5;
  assign rf_matrix_c_1_tile_v_2_MPORT_15_data = rf[rf_matrix_c_1_tile_v_2_MPORT_15_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_1_tile_v_1_MPORT_15_en = handshaked & _GEN_1469;
  assign rf_matrix_c_1_tile_v_1_MPORT_15_addr = 8'ha9;
  assign rf_matrix_c_1_tile_v_1_MPORT_15_data = rf[rf_matrix_c_1_tile_v_1_MPORT_15_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_1_tile_v_0_MPORT_15_en = handshaked & _GEN_1469;
  assign rf_matrix_c_1_tile_v_0_MPORT_15_addr = 8'had;
  assign rf_matrix_c_1_tile_v_0_MPORT_15_data = rf[rf_matrix_c_1_tile_v_0_MPORT_15_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_1_MPORT_40_en = handshaked & _GEN_1483;
  assign rf_a_tile_v_1_MPORT_40_addr = 8'h22;
  assign rf_a_tile_v_1_MPORT_40_data = rf[rf_a_tile_v_1_MPORT_40_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_0_MPORT_40_en = handshaked & _GEN_1483;
  assign rf_a_tile_v_0_MPORT_40_addr = 8'h26;
  assign rf_a_tile_v_0_MPORT_40_data = rf[rf_a_tile_v_0_MPORT_40_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_1_tile_v_3_MPORT_16_en = handshaked & _GEN_1483;
  assign rf_matrix_b_1_tile_v_3_MPORT_16_addr = 8'h60;
  assign rf_matrix_b_1_tile_v_3_MPORT_16_data = rf[rf_matrix_b_1_tile_v_3_MPORT_16_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_1_tile_v_2_MPORT_16_en = handshaked & _GEN_1483;
  assign rf_matrix_b_1_tile_v_2_MPORT_16_addr = 8'h64;
  assign rf_matrix_b_1_tile_v_2_MPORT_16_data = rf[rf_matrix_b_1_tile_v_2_MPORT_16_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_1_tile_v_1_MPORT_16_en = handshaked & _GEN_1483;
  assign rf_matrix_b_1_tile_v_1_MPORT_16_addr = 8'h68;
  assign rf_matrix_b_1_tile_v_1_MPORT_16_data = rf[rf_matrix_b_1_tile_v_1_MPORT_16_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_1_tile_v_0_MPORT_16_en = handshaked & _GEN_1483;
  assign rf_matrix_b_1_tile_v_0_MPORT_16_addr = 8'h6c;
  assign rf_matrix_b_1_tile_v_0_MPORT_16_data = rf[rf_matrix_b_1_tile_v_0_MPORT_16_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_1_tile_v_3_MPORT_16_en = handshaked & _GEN_1483;
  assign rf_matrix_c_1_tile_v_3_MPORT_16_addr = 8'hc2;
  assign rf_matrix_c_1_tile_v_3_MPORT_16_data = rf[rf_matrix_c_1_tile_v_3_MPORT_16_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_1_tile_v_2_MPORT_16_en = handshaked & _GEN_1483;
  assign rf_matrix_c_1_tile_v_2_MPORT_16_addr = 8'hc3;
  assign rf_matrix_c_1_tile_v_2_MPORT_16_data = rf[rf_matrix_c_1_tile_v_2_MPORT_16_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_1_tile_v_1_MPORT_16_en = handshaked & _GEN_1483;
  assign rf_matrix_c_1_tile_v_1_MPORT_16_addr = 8'hca;
  assign rf_matrix_c_1_tile_v_1_MPORT_16_data = rf[rf_matrix_c_1_tile_v_1_MPORT_16_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_1_tile_v_0_MPORT_16_en = handshaked & _GEN_1483;
  assign rf_matrix_c_1_tile_v_0_MPORT_16_addr = 8'hcb;
  assign rf_matrix_c_1_tile_v_0_MPORT_16_data = rf[rf_matrix_c_1_tile_v_0_MPORT_16_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_1_MPORT_41_en = handshaked & _GEN_1495;
  assign rf_a_tile_v_1_MPORT_41_addr = 8'h2a;
  assign rf_a_tile_v_1_MPORT_41_data = rf[rf_a_tile_v_1_MPORT_41_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_0_MPORT_41_en = handshaked & _GEN_1495;
  assign rf_a_tile_v_0_MPORT_41_addr = 8'h2e;
  assign rf_a_tile_v_0_MPORT_41_data = rf[rf_a_tile_v_0_MPORT_41_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_1_tile_v_3_MPORT_17_en = handshaked & _GEN_1495;
  assign rf_matrix_b_1_tile_v_3_MPORT_17_addr = 8'h60;
  assign rf_matrix_b_1_tile_v_3_MPORT_17_data = rf[rf_matrix_b_1_tile_v_3_MPORT_17_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_1_tile_v_2_MPORT_17_en = handshaked & _GEN_1495;
  assign rf_matrix_b_1_tile_v_2_MPORT_17_addr = 8'h64;
  assign rf_matrix_b_1_tile_v_2_MPORT_17_data = rf[rf_matrix_b_1_tile_v_2_MPORT_17_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_1_tile_v_1_MPORT_17_en = handshaked & _GEN_1495;
  assign rf_matrix_b_1_tile_v_1_MPORT_17_addr = 8'h68;
  assign rf_matrix_b_1_tile_v_1_MPORT_17_data = rf[rf_matrix_b_1_tile_v_1_MPORT_17_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_1_tile_v_0_MPORT_17_en = handshaked & _GEN_1495;
  assign rf_matrix_b_1_tile_v_0_MPORT_17_addr = 8'h6c;
  assign rf_matrix_b_1_tile_v_0_MPORT_17_data = rf[rf_matrix_b_1_tile_v_0_MPORT_17_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_1_tile_v_3_MPORT_17_en = handshaked & _GEN_1495;
  assign rf_matrix_c_1_tile_v_3_MPORT_17_addr = 8'hd2;
  assign rf_matrix_c_1_tile_v_3_MPORT_17_data = rf[rf_matrix_c_1_tile_v_3_MPORT_17_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_1_tile_v_2_MPORT_17_en = handshaked & _GEN_1495;
  assign rf_matrix_c_1_tile_v_2_MPORT_17_addr = 8'hd3;
  assign rf_matrix_c_1_tile_v_2_MPORT_17_data = rf[rf_matrix_c_1_tile_v_2_MPORT_17_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_1_tile_v_1_MPORT_17_en = handshaked & _GEN_1495;
  assign rf_matrix_c_1_tile_v_1_MPORT_17_addr = 8'hda;
  assign rf_matrix_c_1_tile_v_1_MPORT_17_data = rf[rf_matrix_c_1_tile_v_1_MPORT_17_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_1_tile_v_0_MPORT_17_en = handshaked & _GEN_1495;
  assign rf_matrix_c_1_tile_v_0_MPORT_17_addr = 8'hdb;
  assign rf_matrix_c_1_tile_v_0_MPORT_17_data = rf[rf_matrix_c_1_tile_v_0_MPORT_17_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_1_MPORT_42_en = handshaked & _GEN_1507;
  assign rf_a_tile_v_1_MPORT_42_addr = 8'h23;
  assign rf_a_tile_v_1_MPORT_42_data = rf[rf_a_tile_v_1_MPORT_42_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_0_MPORT_42_en = handshaked & _GEN_1507;
  assign rf_a_tile_v_0_MPORT_42_addr = 8'h27;
  assign rf_a_tile_v_0_MPORT_42_data = rf[rf_a_tile_v_0_MPORT_42_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_1_tile_v_3_MPORT_18_en = handshaked & _GEN_1507;
  assign rf_matrix_b_1_tile_v_3_MPORT_18_addr = 8'h70;
  assign rf_matrix_b_1_tile_v_3_MPORT_18_data = rf[rf_matrix_b_1_tile_v_3_MPORT_18_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_1_tile_v_2_MPORT_18_en = handshaked & _GEN_1507;
  assign rf_matrix_b_1_tile_v_2_MPORT_18_addr = 8'h74;
  assign rf_matrix_b_1_tile_v_2_MPORT_18_data = rf[rf_matrix_b_1_tile_v_2_MPORT_18_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_1_tile_v_1_MPORT_18_en = handshaked & _GEN_1507;
  assign rf_matrix_b_1_tile_v_1_MPORT_18_addr = 8'h78;
  assign rf_matrix_b_1_tile_v_1_MPORT_18_data = rf[rf_matrix_b_1_tile_v_1_MPORT_18_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_1_tile_v_0_MPORT_18_en = handshaked & _GEN_1507;
  assign rf_matrix_b_1_tile_v_0_MPORT_18_addr = 8'h7c;
  assign rf_matrix_b_1_tile_v_0_MPORT_18_data = rf[rf_matrix_b_1_tile_v_0_MPORT_18_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_1_tile_v_3_MPORT_18_en = handshaked & _GEN_1507;
  assign rf_matrix_c_1_tile_v_3_MPORT_18_addr = 8'hc0;
  assign rf_matrix_c_1_tile_v_3_MPORT_18_data = rf[rf_matrix_c_1_tile_v_3_MPORT_18_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_1_tile_v_2_MPORT_18_en = handshaked & _GEN_1507;
  assign rf_matrix_c_1_tile_v_2_MPORT_18_addr = 8'hc1;
  assign rf_matrix_c_1_tile_v_2_MPORT_18_data = rf[rf_matrix_c_1_tile_v_2_MPORT_18_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_1_tile_v_1_MPORT_18_en = handshaked & _GEN_1507;
  assign rf_matrix_c_1_tile_v_1_MPORT_18_addr = 8'hc8;
  assign rf_matrix_c_1_tile_v_1_MPORT_18_data = rf[rf_matrix_c_1_tile_v_1_MPORT_18_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_1_tile_v_0_MPORT_18_en = handshaked & _GEN_1507;
  assign rf_matrix_c_1_tile_v_0_MPORT_18_addr = 8'hc9;
  assign rf_matrix_c_1_tile_v_0_MPORT_18_data = rf[rf_matrix_c_1_tile_v_0_MPORT_18_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_3_MPORT_14_en = handshaked & _GEN_1519;
  assign rf_a_tile_v_3_MPORT_14_addr = 8'h23;
  assign rf_a_tile_v_3_MPORT_14_data = rf[rf_a_tile_v_3_MPORT_14_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_2_MPORT_14_en = handshaked & _GEN_1519;
  assign rf_a_tile_v_2_MPORT_14_addr = 8'h27;
  assign rf_a_tile_v_2_MPORT_14_data = rf[rf_a_tile_v_2_MPORT_14_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_1_MPORT_43_en = handshaked & _GEN_1519;
  assign rf_a_tile_v_1_MPORT_43_addr = 8'h2b;
  assign rf_a_tile_v_1_MPORT_43_data = rf[rf_a_tile_v_1_MPORT_43_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_0_MPORT_43_en = handshaked & _GEN_1519;
  assign rf_a_tile_v_0_MPORT_43_addr = 8'h2f;
  assign rf_a_tile_v_0_MPORT_43_data = rf[rf_a_tile_v_0_MPORT_43_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_1_tile_v_3_MPORT_19_en = handshaked & _GEN_1519;
  assign rf_matrix_b_1_tile_v_3_MPORT_19_addr = 8'h70;
  assign rf_matrix_b_1_tile_v_3_MPORT_19_data = rf[rf_matrix_b_1_tile_v_3_MPORT_19_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_1_tile_v_2_MPORT_19_en = handshaked & _GEN_1519;
  assign rf_matrix_b_1_tile_v_2_MPORT_19_addr = 8'h74;
  assign rf_matrix_b_1_tile_v_2_MPORT_19_data = rf[rf_matrix_b_1_tile_v_2_MPORT_19_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_1_tile_v_1_MPORT_19_en = handshaked & _GEN_1519;
  assign rf_matrix_b_1_tile_v_1_MPORT_19_addr = 8'h78;
  assign rf_matrix_b_1_tile_v_1_MPORT_19_data = rf[rf_matrix_b_1_tile_v_1_MPORT_19_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_1_tile_v_0_MPORT_19_en = handshaked & _GEN_1519;
  assign rf_matrix_b_1_tile_v_0_MPORT_19_addr = 8'h7c;
  assign rf_matrix_b_1_tile_v_0_MPORT_19_data = rf[rf_matrix_b_1_tile_v_0_MPORT_19_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_1_tile_v_3_MPORT_19_en = handshaked & _GEN_1519;
  assign rf_matrix_c_1_tile_v_3_MPORT_19_addr = 8'ha0;
  assign rf_matrix_c_1_tile_v_3_MPORT_19_data = rf[rf_matrix_c_1_tile_v_3_MPORT_19_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_1_tile_v_2_MPORT_19_en = handshaked & _GEN_1519;
  assign rf_matrix_c_1_tile_v_2_MPORT_19_addr = 8'ha4;
  assign rf_matrix_c_1_tile_v_2_MPORT_19_data = rf[rf_matrix_c_1_tile_v_2_MPORT_19_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_1_tile_v_1_MPORT_19_en = handshaked & _GEN_1519;
  assign rf_matrix_c_1_tile_v_1_MPORT_19_addr = 8'ha8;
  assign rf_matrix_c_1_tile_v_1_MPORT_19_data = rf[rf_matrix_c_1_tile_v_1_MPORT_19_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_1_tile_v_0_MPORT_19_en = handshaked & _GEN_1519;
  assign rf_matrix_c_1_tile_v_0_MPORT_19_addr = 8'hac;
  assign rf_matrix_c_1_tile_v_0_MPORT_19_data = rf[rf_matrix_c_1_tile_v_0_MPORT_19_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_1_MPORT_44_en = handshaked & _GEN_1533;
  assign rf_a_tile_v_1_MPORT_44_addr = 8'h2b;
  assign rf_a_tile_v_1_MPORT_44_data = rf[rf_a_tile_v_1_MPORT_44_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_0_MPORT_44_en = handshaked & _GEN_1533;
  assign rf_a_tile_v_0_MPORT_44_addr = 8'h2f;
  assign rf_a_tile_v_0_MPORT_44_data = rf[rf_a_tile_v_0_MPORT_44_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_1_tile_v_3_MPORT_20_en = handshaked & _GEN_1533;
  assign rf_matrix_b_1_tile_v_3_MPORT_20_addr = 8'h70;
  assign rf_matrix_b_1_tile_v_3_MPORT_20_data = rf[rf_matrix_b_1_tile_v_3_MPORT_20_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_1_tile_v_2_MPORT_20_en = handshaked & _GEN_1533;
  assign rf_matrix_b_1_tile_v_2_MPORT_20_addr = 8'h74;
  assign rf_matrix_b_1_tile_v_2_MPORT_20_data = rf[rf_matrix_b_1_tile_v_2_MPORT_20_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_1_tile_v_1_MPORT_20_en = handshaked & _GEN_1533;
  assign rf_matrix_b_1_tile_v_1_MPORT_20_addr = 8'h78;
  assign rf_matrix_b_1_tile_v_1_MPORT_20_data = rf[rf_matrix_b_1_tile_v_1_MPORT_20_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_1_tile_v_0_MPORT_20_en = handshaked & _GEN_1533;
  assign rf_matrix_b_1_tile_v_0_MPORT_20_addr = 8'h7c;
  assign rf_matrix_b_1_tile_v_0_MPORT_20_data = rf[rf_matrix_b_1_tile_v_0_MPORT_20_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_1_tile_v_3_MPORT_20_en = handshaked & _GEN_1533;
  assign rf_matrix_c_1_tile_v_3_MPORT_20_addr = 8'hd0;
  assign rf_matrix_c_1_tile_v_3_MPORT_20_data = rf[rf_matrix_c_1_tile_v_3_MPORT_20_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_1_tile_v_2_MPORT_20_en = handshaked & _GEN_1533;
  assign rf_matrix_c_1_tile_v_2_MPORT_20_addr = 8'hd1;
  assign rf_matrix_c_1_tile_v_2_MPORT_20_data = rf[rf_matrix_c_1_tile_v_2_MPORT_20_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_1_tile_v_1_MPORT_20_en = handshaked & _GEN_1533;
  assign rf_matrix_c_1_tile_v_1_MPORT_20_addr = 8'hd8;
  assign rf_matrix_c_1_tile_v_1_MPORT_20_data = rf[rf_matrix_c_1_tile_v_1_MPORT_20_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_1_tile_v_0_MPORT_20_en = handshaked & _GEN_1533;
  assign rf_matrix_c_1_tile_v_0_MPORT_20_addr = 8'hd9;
  assign rf_matrix_c_1_tile_v_0_MPORT_20_data = rf[rf_matrix_c_1_tile_v_0_MPORT_20_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_3_MPORT_15_en = handshaked & _GEN_1545;
  assign rf_a_tile_v_3_MPORT_15_addr = 8'h23;
  assign rf_a_tile_v_3_MPORT_15_data = rf[rf_a_tile_v_3_MPORT_15_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_2_MPORT_15_en = handshaked & _GEN_1545;
  assign rf_a_tile_v_2_MPORT_15_addr = 8'h27;
  assign rf_a_tile_v_2_MPORT_15_data = rf[rf_a_tile_v_2_MPORT_15_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_1_MPORT_45_en = handshaked & _GEN_1545;
  assign rf_a_tile_v_1_MPORT_45_addr = 8'h2b;
  assign rf_a_tile_v_1_MPORT_45_data = rf[rf_a_tile_v_1_MPORT_45_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_0_MPORT_45_en = handshaked & _GEN_1545;
  assign rf_a_tile_v_0_MPORT_45_addr = 8'h2f;
  assign rf_a_tile_v_0_MPORT_45_data = rf[rf_a_tile_v_0_MPORT_45_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_1_tile_v_3_MPORT_21_en = handshaked & _GEN_1545;
  assign rf_matrix_b_1_tile_v_3_MPORT_21_addr = 8'h70;
  assign rf_matrix_b_1_tile_v_3_MPORT_21_data = rf[rf_matrix_b_1_tile_v_3_MPORT_21_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_1_tile_v_2_MPORT_21_en = handshaked & _GEN_1545;
  assign rf_matrix_b_1_tile_v_2_MPORT_21_addr = 8'h74;
  assign rf_matrix_b_1_tile_v_2_MPORT_21_data = rf[rf_matrix_b_1_tile_v_2_MPORT_21_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_1_tile_v_1_MPORT_21_en = handshaked & _GEN_1545;
  assign rf_matrix_b_1_tile_v_1_MPORT_21_addr = 8'h78;
  assign rf_matrix_b_1_tile_v_1_MPORT_21_data = rf[rf_matrix_b_1_tile_v_1_MPORT_21_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_1_tile_v_0_MPORT_21_en = handshaked & _GEN_1545;
  assign rf_matrix_b_1_tile_v_0_MPORT_21_addr = 8'h7c;
  assign rf_matrix_b_1_tile_v_0_MPORT_21_data = rf[rf_matrix_b_1_tile_v_0_MPORT_21_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_1_tile_v_3_MPORT_21_en = handshaked & _GEN_1545;
  assign rf_matrix_c_1_tile_v_3_MPORT_21_addr = 8'ha1;
  assign rf_matrix_c_1_tile_v_3_MPORT_21_data = rf[rf_matrix_c_1_tile_v_3_MPORT_21_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_1_tile_v_2_MPORT_21_en = handshaked & _GEN_1545;
  assign rf_matrix_c_1_tile_v_2_MPORT_21_addr = 8'ha5;
  assign rf_matrix_c_1_tile_v_2_MPORT_21_data = rf[rf_matrix_c_1_tile_v_2_MPORT_21_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_1_tile_v_1_MPORT_21_en = handshaked & _GEN_1545;
  assign rf_matrix_c_1_tile_v_1_MPORT_21_addr = 8'ha9;
  assign rf_matrix_c_1_tile_v_1_MPORT_21_data = rf[rf_matrix_c_1_tile_v_1_MPORT_21_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_1_tile_v_0_MPORT_21_en = handshaked & _GEN_1545;
  assign rf_matrix_c_1_tile_v_0_MPORT_21_addr = 8'had;
  assign rf_matrix_c_1_tile_v_0_MPORT_21_data = rf[rf_matrix_c_1_tile_v_0_MPORT_21_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_1_MPORT_46_en = handshaked & _GEN_1559;
  assign rf_a_tile_v_1_MPORT_46_addr = 8'h23;
  assign rf_a_tile_v_1_MPORT_46_data = rf[rf_a_tile_v_1_MPORT_46_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_0_MPORT_46_en = handshaked & _GEN_1559;
  assign rf_a_tile_v_0_MPORT_46_addr = 8'h27;
  assign rf_a_tile_v_0_MPORT_46_data = rf[rf_a_tile_v_0_MPORT_46_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_1_tile_v_3_MPORT_22_en = handshaked & _GEN_1559;
  assign rf_matrix_b_1_tile_v_3_MPORT_22_addr = 8'h70;
  assign rf_matrix_b_1_tile_v_3_MPORT_22_data = rf[rf_matrix_b_1_tile_v_3_MPORT_22_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_1_tile_v_2_MPORT_22_en = handshaked & _GEN_1559;
  assign rf_matrix_b_1_tile_v_2_MPORT_22_addr = 8'h74;
  assign rf_matrix_b_1_tile_v_2_MPORT_22_data = rf[rf_matrix_b_1_tile_v_2_MPORT_22_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_1_tile_v_1_MPORT_22_en = handshaked & _GEN_1559;
  assign rf_matrix_b_1_tile_v_1_MPORT_22_addr = 8'h78;
  assign rf_matrix_b_1_tile_v_1_MPORT_22_data = rf[rf_matrix_b_1_tile_v_1_MPORT_22_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_1_tile_v_0_MPORT_22_en = handshaked & _GEN_1559;
  assign rf_matrix_b_1_tile_v_0_MPORT_22_addr = 8'h7c;
  assign rf_matrix_b_1_tile_v_0_MPORT_22_data = rf[rf_matrix_b_1_tile_v_0_MPORT_22_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_1_tile_v_3_MPORT_22_en = handshaked & _GEN_1559;
  assign rf_matrix_c_1_tile_v_3_MPORT_22_addr = 8'hc2;
  assign rf_matrix_c_1_tile_v_3_MPORT_22_data = rf[rf_matrix_c_1_tile_v_3_MPORT_22_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_1_tile_v_2_MPORT_22_en = handshaked & _GEN_1559;
  assign rf_matrix_c_1_tile_v_2_MPORT_22_addr = 8'hc3;
  assign rf_matrix_c_1_tile_v_2_MPORT_22_data = rf[rf_matrix_c_1_tile_v_2_MPORT_22_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_1_tile_v_1_MPORT_22_en = handshaked & _GEN_1559;
  assign rf_matrix_c_1_tile_v_1_MPORT_22_addr = 8'hca;
  assign rf_matrix_c_1_tile_v_1_MPORT_22_data = rf[rf_matrix_c_1_tile_v_1_MPORT_22_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_1_tile_v_0_MPORT_22_en = handshaked & _GEN_1559;
  assign rf_matrix_c_1_tile_v_0_MPORT_22_addr = 8'hcb;
  assign rf_matrix_c_1_tile_v_0_MPORT_22_data = rf[rf_matrix_c_1_tile_v_0_MPORT_22_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_1_MPORT_47_en = handshaked & _GEN_1571;
  assign rf_a_tile_v_1_MPORT_47_addr = 8'h2b;
  assign rf_a_tile_v_1_MPORT_47_data = rf[rf_a_tile_v_1_MPORT_47_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_0_MPORT_47_en = handshaked & _GEN_1571;
  assign rf_a_tile_v_0_MPORT_47_addr = 8'h2f;
  assign rf_a_tile_v_0_MPORT_47_data = rf[rf_a_tile_v_0_MPORT_47_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_1_tile_v_3_MPORT_23_en = handshaked & _GEN_1571;
  assign rf_matrix_b_1_tile_v_3_MPORT_23_addr = 8'h70;
  assign rf_matrix_b_1_tile_v_3_MPORT_23_data = rf[rf_matrix_b_1_tile_v_3_MPORT_23_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_1_tile_v_2_MPORT_23_en = handshaked & _GEN_1571;
  assign rf_matrix_b_1_tile_v_2_MPORT_23_addr = 8'h74;
  assign rf_matrix_b_1_tile_v_2_MPORT_23_data = rf[rf_matrix_b_1_tile_v_2_MPORT_23_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_1_tile_v_1_MPORT_23_en = handshaked & _GEN_1571;
  assign rf_matrix_b_1_tile_v_1_MPORT_23_addr = 8'h78;
  assign rf_matrix_b_1_tile_v_1_MPORT_23_data = rf[rf_matrix_b_1_tile_v_1_MPORT_23_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_1_tile_v_0_MPORT_23_en = handshaked & _GEN_1571;
  assign rf_matrix_b_1_tile_v_0_MPORT_23_addr = 8'h7c;
  assign rf_matrix_b_1_tile_v_0_MPORT_23_data = rf[rf_matrix_b_1_tile_v_0_MPORT_23_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_1_tile_v_3_MPORT_23_en = handshaked & _GEN_1571;
  assign rf_matrix_c_1_tile_v_3_MPORT_23_addr = 8'hd2;
  assign rf_matrix_c_1_tile_v_3_MPORT_23_data = rf[rf_matrix_c_1_tile_v_3_MPORT_23_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_1_tile_v_2_MPORT_23_en = handshaked & _GEN_1571;
  assign rf_matrix_c_1_tile_v_2_MPORT_23_addr = 8'hd3;
  assign rf_matrix_c_1_tile_v_2_MPORT_23_data = rf[rf_matrix_c_1_tile_v_2_MPORT_23_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_1_tile_v_1_MPORT_23_en = handshaked & _GEN_1571;
  assign rf_matrix_c_1_tile_v_1_MPORT_23_addr = 8'hda;
  assign rf_matrix_c_1_tile_v_1_MPORT_23_data = rf[rf_matrix_c_1_tile_v_1_MPORT_23_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_1_tile_v_0_MPORT_23_en = handshaked & _GEN_1571;
  assign rf_matrix_c_1_tile_v_0_MPORT_23_addr = 8'hdb;
  assign rf_matrix_c_1_tile_v_0_MPORT_23_data = rf[rf_matrix_c_1_tile_v_0_MPORT_23_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_1_MPORT_48_en = handshaked & _GEN_1276;
  assign rf_a_tile_v_1_MPORT_48_addr = 8'h0;
  assign rf_a_tile_v_1_MPORT_48_data = rf[rf_a_tile_v_1_MPORT_48_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_0_MPORT_48_en = handshaked & _GEN_1276;
  assign rf_a_tile_v_0_MPORT_48_addr = 8'h4;
  assign rf_a_tile_v_0_MPORT_48_data = rf[rf_a_tile_v_0_MPORT_48_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_2_tile_v_3_MPORT_en = handshaked & _GEN_1276;
  assign rf_matrix_b_2_tile_v_3_MPORT_addr = 8'h42;
  assign rf_matrix_b_2_tile_v_3_MPORT_data = rf[rf_matrix_b_2_tile_v_3_MPORT_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_2_tile_v_2_MPORT_en = handshaked & _GEN_1276;
  assign rf_matrix_b_2_tile_v_2_MPORT_addr = 8'h46;
  assign rf_matrix_b_2_tile_v_2_MPORT_data = rf[rf_matrix_b_2_tile_v_2_MPORT_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_2_tile_v_1_MPORT_en = handshaked & _GEN_1276;
  assign rf_matrix_b_2_tile_v_1_MPORT_addr = 8'h4a;
  assign rf_matrix_b_2_tile_v_1_MPORT_data = rf[rf_matrix_b_2_tile_v_1_MPORT_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_2_tile_v_0_MPORT_en = handshaked & _GEN_1276;
  assign rf_matrix_b_2_tile_v_0_MPORT_addr = 8'h4e;
  assign rf_matrix_b_2_tile_v_0_MPORT_data = rf[rf_matrix_b_2_tile_v_0_MPORT_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_2_tile_v_3_MPORT_en = handshaked & _GEN_1276;
  assign rf_matrix_c_2_tile_v_3_MPORT_addr = 8'h84;
  assign rf_matrix_c_2_tile_v_3_MPORT_data = rf[rf_matrix_c_2_tile_v_3_MPORT_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_2_tile_v_2_MPORT_en = handshaked & _GEN_1276;
  assign rf_matrix_c_2_tile_v_2_MPORT_addr = 8'h85;
  assign rf_matrix_c_2_tile_v_2_MPORT_data = rf[rf_matrix_c_2_tile_v_2_MPORT_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_2_tile_v_1_MPORT_en = handshaked & _GEN_1276;
  assign rf_matrix_c_2_tile_v_1_MPORT_addr = 8'h8c;
  assign rf_matrix_c_2_tile_v_1_MPORT_data = rf[rf_matrix_c_2_tile_v_1_MPORT_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_2_tile_v_0_MPORT_en = handshaked & _GEN_1276;
  assign rf_matrix_c_2_tile_v_0_MPORT_addr = 8'h8d;
  assign rf_matrix_c_2_tile_v_0_MPORT_data = rf[rf_matrix_c_2_tile_v_0_MPORT_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_3_MPORT_16_en = handshaked & _GEN_1291;
  assign rf_a_tile_v_3_MPORT_16_addr = 8'h0;
  assign rf_a_tile_v_3_MPORT_16_data = rf[rf_a_tile_v_3_MPORT_16_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_2_MPORT_16_en = handshaked & _GEN_1291;
  assign rf_a_tile_v_2_MPORT_16_addr = 8'h4;
  assign rf_a_tile_v_2_MPORT_16_data = rf[rf_a_tile_v_2_MPORT_16_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_1_MPORT_49_en = handshaked & _GEN_1291;
  assign rf_a_tile_v_1_MPORT_49_addr = 8'h8;
  assign rf_a_tile_v_1_MPORT_49_data = rf[rf_a_tile_v_1_MPORT_49_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_0_MPORT_49_en = handshaked & _GEN_1291;
  assign rf_a_tile_v_0_MPORT_49_addr = 8'hc;
  assign rf_a_tile_v_0_MPORT_49_data = rf[rf_a_tile_v_0_MPORT_49_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_2_tile_v_3_MPORT_1_en = handshaked & _GEN_1291;
  assign rf_matrix_b_2_tile_v_3_MPORT_1_addr = 8'h42;
  assign rf_matrix_b_2_tile_v_3_MPORT_1_data = rf[rf_matrix_b_2_tile_v_3_MPORT_1_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_2_tile_v_2_MPORT_1_en = handshaked & _GEN_1291;
  assign rf_matrix_b_2_tile_v_2_MPORT_1_addr = 8'h46;
  assign rf_matrix_b_2_tile_v_2_MPORT_1_data = rf[rf_matrix_b_2_tile_v_2_MPORT_1_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_2_tile_v_1_MPORT_1_en = handshaked & _GEN_1291;
  assign rf_matrix_b_2_tile_v_1_MPORT_1_addr = 8'h4a;
  assign rf_matrix_b_2_tile_v_1_MPORT_1_data = rf[rf_matrix_b_2_tile_v_1_MPORT_1_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_2_tile_v_0_MPORT_1_en = handshaked & _GEN_1291;
  assign rf_matrix_b_2_tile_v_0_MPORT_1_addr = 8'h4e;
  assign rf_matrix_b_2_tile_v_0_MPORT_1_data = rf[rf_matrix_b_2_tile_v_0_MPORT_1_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_2_tile_v_3_MPORT_1_en = handshaked & _GEN_1291;
  assign rf_matrix_c_2_tile_v_3_MPORT_1_addr = 8'h82;
  assign rf_matrix_c_2_tile_v_3_MPORT_1_data = rf[rf_matrix_c_2_tile_v_3_MPORT_1_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_2_tile_v_2_MPORT_1_en = handshaked & _GEN_1291;
  assign rf_matrix_c_2_tile_v_2_MPORT_1_addr = 8'h86;
  assign rf_matrix_c_2_tile_v_2_MPORT_1_data = rf[rf_matrix_c_2_tile_v_2_MPORT_1_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_2_tile_v_1_MPORT_1_en = handshaked & _GEN_1291;
  assign rf_matrix_c_2_tile_v_1_MPORT_1_addr = 8'h8a;
  assign rf_matrix_c_2_tile_v_1_MPORT_1_data = rf[rf_matrix_c_2_tile_v_1_MPORT_1_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_2_tile_v_0_MPORT_1_en = handshaked & _GEN_1291;
  assign rf_matrix_c_2_tile_v_0_MPORT_1_addr = 8'h8e;
  assign rf_matrix_c_2_tile_v_0_MPORT_1_data = rf[rf_matrix_c_2_tile_v_0_MPORT_1_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_1_MPORT_50_en = handshaked & _GEN_1305;
  assign rf_a_tile_v_1_MPORT_50_addr = 8'h8;
  assign rf_a_tile_v_1_MPORT_50_data = rf[rf_a_tile_v_1_MPORT_50_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_0_MPORT_50_en = handshaked & _GEN_1305;
  assign rf_a_tile_v_0_MPORT_50_addr = 8'hc;
  assign rf_a_tile_v_0_MPORT_50_data = rf[rf_a_tile_v_0_MPORT_50_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_2_tile_v_3_MPORT_2_en = handshaked & _GEN_1305;
  assign rf_matrix_b_2_tile_v_3_MPORT_2_addr = 8'h42;
  assign rf_matrix_b_2_tile_v_3_MPORT_2_data = rf[rf_matrix_b_2_tile_v_3_MPORT_2_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_2_tile_v_2_MPORT_2_en = handshaked & _GEN_1305;
  assign rf_matrix_b_2_tile_v_2_MPORT_2_addr = 8'h46;
  assign rf_matrix_b_2_tile_v_2_MPORT_2_data = rf[rf_matrix_b_2_tile_v_2_MPORT_2_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_2_tile_v_1_MPORT_2_en = handshaked & _GEN_1305;
  assign rf_matrix_b_2_tile_v_1_MPORT_2_addr = 8'h4a;
  assign rf_matrix_b_2_tile_v_1_MPORT_2_data = rf[rf_matrix_b_2_tile_v_1_MPORT_2_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_2_tile_v_0_MPORT_2_en = handshaked & _GEN_1305;
  assign rf_matrix_b_2_tile_v_0_MPORT_2_addr = 8'h4e;
  assign rf_matrix_b_2_tile_v_0_MPORT_2_data = rf[rf_matrix_b_2_tile_v_0_MPORT_2_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_2_tile_v_3_MPORT_2_en = handshaked & _GEN_1305;
  assign rf_matrix_c_2_tile_v_3_MPORT_2_addr = 8'h94;
  assign rf_matrix_c_2_tile_v_3_MPORT_2_data = rf[rf_matrix_c_2_tile_v_3_MPORT_2_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_2_tile_v_2_MPORT_2_en = handshaked & _GEN_1305;
  assign rf_matrix_c_2_tile_v_2_MPORT_2_addr = 8'h95;
  assign rf_matrix_c_2_tile_v_2_MPORT_2_data = rf[rf_matrix_c_2_tile_v_2_MPORT_2_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_2_tile_v_1_MPORT_2_en = handshaked & _GEN_1305;
  assign rf_matrix_c_2_tile_v_1_MPORT_2_addr = 8'h9c;
  assign rf_matrix_c_2_tile_v_1_MPORT_2_data = rf[rf_matrix_c_2_tile_v_1_MPORT_2_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_2_tile_v_0_MPORT_2_en = handshaked & _GEN_1305;
  assign rf_matrix_c_2_tile_v_0_MPORT_2_addr = 8'h9d;
  assign rf_matrix_c_2_tile_v_0_MPORT_2_data = rf[rf_matrix_c_2_tile_v_0_MPORT_2_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_3_MPORT_17_en = handshaked & _GEN_1317;
  assign rf_a_tile_v_3_MPORT_17_addr = 8'h0;
  assign rf_a_tile_v_3_MPORT_17_data = rf[rf_a_tile_v_3_MPORT_17_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_2_MPORT_17_en = handshaked & _GEN_1317;
  assign rf_a_tile_v_2_MPORT_17_addr = 8'h4;
  assign rf_a_tile_v_2_MPORT_17_data = rf[rf_a_tile_v_2_MPORT_17_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_1_MPORT_51_en = handshaked & _GEN_1317;
  assign rf_a_tile_v_1_MPORT_51_addr = 8'h8;
  assign rf_a_tile_v_1_MPORT_51_data = rf[rf_a_tile_v_1_MPORT_51_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_0_MPORT_51_en = handshaked & _GEN_1317;
  assign rf_a_tile_v_0_MPORT_51_addr = 8'hc;
  assign rf_a_tile_v_0_MPORT_51_data = rf[rf_a_tile_v_0_MPORT_51_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_2_tile_v_3_MPORT_3_en = handshaked & _GEN_1317;
  assign rf_matrix_b_2_tile_v_3_MPORT_3_addr = 8'h42;
  assign rf_matrix_b_2_tile_v_3_MPORT_3_data = rf[rf_matrix_b_2_tile_v_3_MPORT_3_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_2_tile_v_2_MPORT_3_en = handshaked & _GEN_1317;
  assign rf_matrix_b_2_tile_v_2_MPORT_3_addr = 8'h46;
  assign rf_matrix_b_2_tile_v_2_MPORT_3_data = rf[rf_matrix_b_2_tile_v_2_MPORT_3_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_2_tile_v_1_MPORT_3_en = handshaked & _GEN_1317;
  assign rf_matrix_b_2_tile_v_1_MPORT_3_addr = 8'h4a;
  assign rf_matrix_b_2_tile_v_1_MPORT_3_data = rf[rf_matrix_b_2_tile_v_1_MPORT_3_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_2_tile_v_0_MPORT_3_en = handshaked & _GEN_1317;
  assign rf_matrix_b_2_tile_v_0_MPORT_3_addr = 8'h4e;
  assign rf_matrix_b_2_tile_v_0_MPORT_3_data = rf[rf_matrix_b_2_tile_v_0_MPORT_3_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_2_tile_v_3_MPORT_3_en = handshaked & _GEN_1317;
  assign rf_matrix_c_2_tile_v_3_MPORT_3_addr = 8'h83;
  assign rf_matrix_c_2_tile_v_3_MPORT_3_data = rf[rf_matrix_c_2_tile_v_3_MPORT_3_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_2_tile_v_2_MPORT_3_en = handshaked & _GEN_1317;
  assign rf_matrix_c_2_tile_v_2_MPORT_3_addr = 8'h87;
  assign rf_matrix_c_2_tile_v_2_MPORT_3_data = rf[rf_matrix_c_2_tile_v_2_MPORT_3_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_2_tile_v_1_MPORT_3_en = handshaked & _GEN_1317;
  assign rf_matrix_c_2_tile_v_1_MPORT_3_addr = 8'h8b;
  assign rf_matrix_c_2_tile_v_1_MPORT_3_data = rf[rf_matrix_c_2_tile_v_1_MPORT_3_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_2_tile_v_0_MPORT_3_en = handshaked & _GEN_1317;
  assign rf_matrix_c_2_tile_v_0_MPORT_3_addr = 8'h8f;
  assign rf_matrix_c_2_tile_v_0_MPORT_3_data = rf[rf_matrix_c_2_tile_v_0_MPORT_3_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_1_MPORT_52_en = handshaked & _GEN_1331;
  assign rf_a_tile_v_1_MPORT_52_addr = 8'h0;
  assign rf_a_tile_v_1_MPORT_52_data = rf[rf_a_tile_v_1_MPORT_52_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_0_MPORT_52_en = handshaked & _GEN_1331;
  assign rf_a_tile_v_0_MPORT_52_addr = 8'h4;
  assign rf_a_tile_v_0_MPORT_52_data = rf[rf_a_tile_v_0_MPORT_52_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_2_tile_v_3_MPORT_4_en = handshaked & _GEN_1331;
  assign rf_matrix_b_2_tile_v_3_MPORT_4_addr = 8'h42;
  assign rf_matrix_b_2_tile_v_3_MPORT_4_data = rf[rf_matrix_b_2_tile_v_3_MPORT_4_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_2_tile_v_2_MPORT_4_en = handshaked & _GEN_1331;
  assign rf_matrix_b_2_tile_v_2_MPORT_4_addr = 8'h46;
  assign rf_matrix_b_2_tile_v_2_MPORT_4_data = rf[rf_matrix_b_2_tile_v_2_MPORT_4_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_2_tile_v_1_MPORT_4_en = handshaked & _GEN_1331;
  assign rf_matrix_b_2_tile_v_1_MPORT_4_addr = 8'h4a;
  assign rf_matrix_b_2_tile_v_1_MPORT_4_data = rf[rf_matrix_b_2_tile_v_1_MPORT_4_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_2_tile_v_0_MPORT_4_en = handshaked & _GEN_1331;
  assign rf_matrix_b_2_tile_v_0_MPORT_4_addr = 8'h4e;
  assign rf_matrix_b_2_tile_v_0_MPORT_4_data = rf[rf_matrix_b_2_tile_v_0_MPORT_4_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_2_tile_v_3_MPORT_4_en = handshaked & _GEN_1331;
  assign rf_matrix_c_2_tile_v_3_MPORT_4_addr = 8'h86;
  assign rf_matrix_c_2_tile_v_3_MPORT_4_data = rf[rf_matrix_c_2_tile_v_3_MPORT_4_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_2_tile_v_2_MPORT_4_en = handshaked & _GEN_1331;
  assign rf_matrix_c_2_tile_v_2_MPORT_4_addr = 8'h87;
  assign rf_matrix_c_2_tile_v_2_MPORT_4_data = rf[rf_matrix_c_2_tile_v_2_MPORT_4_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_2_tile_v_1_MPORT_4_en = handshaked & _GEN_1331;
  assign rf_matrix_c_2_tile_v_1_MPORT_4_addr = 8'h8e;
  assign rf_matrix_c_2_tile_v_1_MPORT_4_data = rf[rf_matrix_c_2_tile_v_1_MPORT_4_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_2_tile_v_0_MPORT_4_en = handshaked & _GEN_1331;
  assign rf_matrix_c_2_tile_v_0_MPORT_4_addr = 8'h8f;
  assign rf_matrix_c_2_tile_v_0_MPORT_4_data = rf[rf_matrix_c_2_tile_v_0_MPORT_4_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_1_MPORT_53_en = handshaked & _GEN_1343;
  assign rf_a_tile_v_1_MPORT_53_addr = 8'h8;
  assign rf_a_tile_v_1_MPORT_53_data = rf[rf_a_tile_v_1_MPORT_53_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_0_MPORT_53_en = handshaked & _GEN_1343;
  assign rf_a_tile_v_0_MPORT_53_addr = 8'hc;
  assign rf_a_tile_v_0_MPORT_53_data = rf[rf_a_tile_v_0_MPORT_53_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_2_tile_v_3_MPORT_5_en = handshaked & _GEN_1343;
  assign rf_matrix_b_2_tile_v_3_MPORT_5_addr = 8'h42;
  assign rf_matrix_b_2_tile_v_3_MPORT_5_data = rf[rf_matrix_b_2_tile_v_3_MPORT_5_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_2_tile_v_2_MPORT_5_en = handshaked & _GEN_1343;
  assign rf_matrix_b_2_tile_v_2_MPORT_5_addr = 8'h46;
  assign rf_matrix_b_2_tile_v_2_MPORT_5_data = rf[rf_matrix_b_2_tile_v_2_MPORT_5_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_2_tile_v_1_MPORT_5_en = handshaked & _GEN_1343;
  assign rf_matrix_b_2_tile_v_1_MPORT_5_addr = 8'h4a;
  assign rf_matrix_b_2_tile_v_1_MPORT_5_data = rf[rf_matrix_b_2_tile_v_1_MPORT_5_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_2_tile_v_0_MPORT_5_en = handshaked & _GEN_1343;
  assign rf_matrix_b_2_tile_v_0_MPORT_5_addr = 8'h4e;
  assign rf_matrix_b_2_tile_v_0_MPORT_5_data = rf[rf_matrix_b_2_tile_v_0_MPORT_5_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_2_tile_v_3_MPORT_5_en = handshaked & _GEN_1343;
  assign rf_matrix_c_2_tile_v_3_MPORT_5_addr = 8'h96;
  assign rf_matrix_c_2_tile_v_3_MPORT_5_data = rf[rf_matrix_c_2_tile_v_3_MPORT_5_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_2_tile_v_2_MPORT_5_en = handshaked & _GEN_1343;
  assign rf_matrix_c_2_tile_v_2_MPORT_5_addr = 8'h97;
  assign rf_matrix_c_2_tile_v_2_MPORT_5_data = rf[rf_matrix_c_2_tile_v_2_MPORT_5_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_2_tile_v_1_MPORT_5_en = handshaked & _GEN_1343;
  assign rf_matrix_c_2_tile_v_1_MPORT_5_addr = 8'h9e;
  assign rf_matrix_c_2_tile_v_1_MPORT_5_data = rf[rf_matrix_c_2_tile_v_1_MPORT_5_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_2_tile_v_0_MPORT_5_en = handshaked & _GEN_1343;
  assign rf_matrix_c_2_tile_v_0_MPORT_5_addr = 8'h9f;
  assign rf_matrix_c_2_tile_v_0_MPORT_5_data = rf[rf_matrix_c_2_tile_v_0_MPORT_5_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_1_MPORT_54_en = handshaked & _GEN_1355;
  assign rf_a_tile_v_1_MPORT_54_addr = 8'h1;
  assign rf_a_tile_v_1_MPORT_54_data = rf[rf_a_tile_v_1_MPORT_54_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_0_MPORT_54_en = handshaked & _GEN_1355;
  assign rf_a_tile_v_0_MPORT_54_addr = 8'h5;
  assign rf_a_tile_v_0_MPORT_54_data = rf[rf_a_tile_v_0_MPORT_54_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_2_tile_v_3_MPORT_6_en = handshaked & _GEN_1355;
  assign rf_matrix_b_2_tile_v_3_MPORT_6_addr = 8'h52;
  assign rf_matrix_b_2_tile_v_3_MPORT_6_data = rf[rf_matrix_b_2_tile_v_3_MPORT_6_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_2_tile_v_2_MPORT_6_en = handshaked & _GEN_1355;
  assign rf_matrix_b_2_tile_v_2_MPORT_6_addr = 8'h56;
  assign rf_matrix_b_2_tile_v_2_MPORT_6_data = rf[rf_matrix_b_2_tile_v_2_MPORT_6_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_2_tile_v_1_MPORT_6_en = handshaked & _GEN_1355;
  assign rf_matrix_b_2_tile_v_1_MPORT_6_addr = 8'h5a;
  assign rf_matrix_b_2_tile_v_1_MPORT_6_data = rf[rf_matrix_b_2_tile_v_1_MPORT_6_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_2_tile_v_0_MPORT_6_en = handshaked & _GEN_1355;
  assign rf_matrix_b_2_tile_v_0_MPORT_6_addr = 8'h5e;
  assign rf_matrix_b_2_tile_v_0_MPORT_6_data = rf[rf_matrix_b_2_tile_v_0_MPORT_6_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_2_tile_v_3_MPORT_6_en = handshaked & _GEN_1355;
  assign rf_matrix_c_2_tile_v_3_MPORT_6_addr = 8'h84;
  assign rf_matrix_c_2_tile_v_3_MPORT_6_data = rf[rf_matrix_c_2_tile_v_3_MPORT_6_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_2_tile_v_2_MPORT_6_en = handshaked & _GEN_1355;
  assign rf_matrix_c_2_tile_v_2_MPORT_6_addr = 8'h85;
  assign rf_matrix_c_2_tile_v_2_MPORT_6_data = rf[rf_matrix_c_2_tile_v_2_MPORT_6_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_2_tile_v_1_MPORT_6_en = handshaked & _GEN_1355;
  assign rf_matrix_c_2_tile_v_1_MPORT_6_addr = 8'h8c;
  assign rf_matrix_c_2_tile_v_1_MPORT_6_data = rf[rf_matrix_c_2_tile_v_1_MPORT_6_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_2_tile_v_0_MPORT_6_en = handshaked & _GEN_1355;
  assign rf_matrix_c_2_tile_v_0_MPORT_6_addr = 8'h8d;
  assign rf_matrix_c_2_tile_v_0_MPORT_6_data = rf[rf_matrix_c_2_tile_v_0_MPORT_6_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_3_MPORT_18_en = handshaked & _GEN_1367;
  assign rf_a_tile_v_3_MPORT_18_addr = 8'h1;
  assign rf_a_tile_v_3_MPORT_18_data = rf[rf_a_tile_v_3_MPORT_18_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_2_MPORT_18_en = handshaked & _GEN_1367;
  assign rf_a_tile_v_2_MPORT_18_addr = 8'h5;
  assign rf_a_tile_v_2_MPORT_18_data = rf[rf_a_tile_v_2_MPORT_18_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_1_MPORT_55_en = handshaked & _GEN_1367;
  assign rf_a_tile_v_1_MPORT_55_addr = 8'h9;
  assign rf_a_tile_v_1_MPORT_55_data = rf[rf_a_tile_v_1_MPORT_55_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_0_MPORT_55_en = handshaked & _GEN_1367;
  assign rf_a_tile_v_0_MPORT_55_addr = 8'hd;
  assign rf_a_tile_v_0_MPORT_55_data = rf[rf_a_tile_v_0_MPORT_55_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_2_tile_v_3_MPORT_7_en = handshaked & _GEN_1367;
  assign rf_matrix_b_2_tile_v_3_MPORT_7_addr = 8'h52;
  assign rf_matrix_b_2_tile_v_3_MPORT_7_data = rf[rf_matrix_b_2_tile_v_3_MPORT_7_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_2_tile_v_2_MPORT_7_en = handshaked & _GEN_1367;
  assign rf_matrix_b_2_tile_v_2_MPORT_7_addr = 8'h56;
  assign rf_matrix_b_2_tile_v_2_MPORT_7_data = rf[rf_matrix_b_2_tile_v_2_MPORT_7_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_2_tile_v_1_MPORT_7_en = handshaked & _GEN_1367;
  assign rf_matrix_b_2_tile_v_1_MPORT_7_addr = 8'h5a;
  assign rf_matrix_b_2_tile_v_1_MPORT_7_data = rf[rf_matrix_b_2_tile_v_1_MPORT_7_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_2_tile_v_0_MPORT_7_en = handshaked & _GEN_1367;
  assign rf_matrix_b_2_tile_v_0_MPORT_7_addr = 8'h5e;
  assign rf_matrix_b_2_tile_v_0_MPORT_7_data = rf[rf_matrix_b_2_tile_v_0_MPORT_7_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_2_tile_v_3_MPORT_7_en = handshaked & _GEN_1367;
  assign rf_matrix_c_2_tile_v_3_MPORT_7_addr = 8'h82;
  assign rf_matrix_c_2_tile_v_3_MPORT_7_data = rf[rf_matrix_c_2_tile_v_3_MPORT_7_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_2_tile_v_2_MPORT_7_en = handshaked & _GEN_1367;
  assign rf_matrix_c_2_tile_v_2_MPORT_7_addr = 8'h86;
  assign rf_matrix_c_2_tile_v_2_MPORT_7_data = rf[rf_matrix_c_2_tile_v_2_MPORT_7_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_2_tile_v_1_MPORT_7_en = handshaked & _GEN_1367;
  assign rf_matrix_c_2_tile_v_1_MPORT_7_addr = 8'h8a;
  assign rf_matrix_c_2_tile_v_1_MPORT_7_data = rf[rf_matrix_c_2_tile_v_1_MPORT_7_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_2_tile_v_0_MPORT_7_en = handshaked & _GEN_1367;
  assign rf_matrix_c_2_tile_v_0_MPORT_7_addr = 8'h8e;
  assign rf_matrix_c_2_tile_v_0_MPORT_7_data = rf[rf_matrix_c_2_tile_v_0_MPORT_7_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_1_MPORT_56_en = handshaked & _GEN_1381;
  assign rf_a_tile_v_1_MPORT_56_addr = 8'h9;
  assign rf_a_tile_v_1_MPORT_56_data = rf[rf_a_tile_v_1_MPORT_56_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_0_MPORT_56_en = handshaked & _GEN_1381;
  assign rf_a_tile_v_0_MPORT_56_addr = 8'hd;
  assign rf_a_tile_v_0_MPORT_56_data = rf[rf_a_tile_v_0_MPORT_56_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_2_tile_v_3_MPORT_8_en = handshaked & _GEN_1381;
  assign rf_matrix_b_2_tile_v_3_MPORT_8_addr = 8'h52;
  assign rf_matrix_b_2_tile_v_3_MPORT_8_data = rf[rf_matrix_b_2_tile_v_3_MPORT_8_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_2_tile_v_2_MPORT_8_en = handshaked & _GEN_1381;
  assign rf_matrix_b_2_tile_v_2_MPORT_8_addr = 8'h56;
  assign rf_matrix_b_2_tile_v_2_MPORT_8_data = rf[rf_matrix_b_2_tile_v_2_MPORT_8_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_2_tile_v_1_MPORT_8_en = handshaked & _GEN_1381;
  assign rf_matrix_b_2_tile_v_1_MPORT_8_addr = 8'h5a;
  assign rf_matrix_b_2_tile_v_1_MPORT_8_data = rf[rf_matrix_b_2_tile_v_1_MPORT_8_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_2_tile_v_0_MPORT_8_en = handshaked & _GEN_1381;
  assign rf_matrix_b_2_tile_v_0_MPORT_8_addr = 8'h5e;
  assign rf_matrix_b_2_tile_v_0_MPORT_8_data = rf[rf_matrix_b_2_tile_v_0_MPORT_8_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_2_tile_v_3_MPORT_8_en = handshaked & _GEN_1381;
  assign rf_matrix_c_2_tile_v_3_MPORT_8_addr = 8'h94;
  assign rf_matrix_c_2_tile_v_3_MPORT_8_data = rf[rf_matrix_c_2_tile_v_3_MPORT_8_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_2_tile_v_2_MPORT_8_en = handshaked & _GEN_1381;
  assign rf_matrix_c_2_tile_v_2_MPORT_8_addr = 8'h95;
  assign rf_matrix_c_2_tile_v_2_MPORT_8_data = rf[rf_matrix_c_2_tile_v_2_MPORT_8_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_2_tile_v_1_MPORT_8_en = handshaked & _GEN_1381;
  assign rf_matrix_c_2_tile_v_1_MPORT_8_addr = 8'h9c;
  assign rf_matrix_c_2_tile_v_1_MPORT_8_data = rf[rf_matrix_c_2_tile_v_1_MPORT_8_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_2_tile_v_0_MPORT_8_en = handshaked & _GEN_1381;
  assign rf_matrix_c_2_tile_v_0_MPORT_8_addr = 8'h9d;
  assign rf_matrix_c_2_tile_v_0_MPORT_8_data = rf[rf_matrix_c_2_tile_v_0_MPORT_8_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_3_MPORT_19_en = handshaked & _GEN_1393;
  assign rf_a_tile_v_3_MPORT_19_addr = 8'h1;
  assign rf_a_tile_v_3_MPORT_19_data = rf[rf_a_tile_v_3_MPORT_19_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_2_MPORT_19_en = handshaked & _GEN_1393;
  assign rf_a_tile_v_2_MPORT_19_addr = 8'h5;
  assign rf_a_tile_v_2_MPORT_19_data = rf[rf_a_tile_v_2_MPORT_19_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_1_MPORT_57_en = handshaked & _GEN_1393;
  assign rf_a_tile_v_1_MPORT_57_addr = 8'h9;
  assign rf_a_tile_v_1_MPORT_57_data = rf[rf_a_tile_v_1_MPORT_57_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_0_MPORT_57_en = handshaked & _GEN_1393;
  assign rf_a_tile_v_0_MPORT_57_addr = 8'hd;
  assign rf_a_tile_v_0_MPORT_57_data = rf[rf_a_tile_v_0_MPORT_57_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_2_tile_v_3_MPORT_9_en = handshaked & _GEN_1393;
  assign rf_matrix_b_2_tile_v_3_MPORT_9_addr = 8'h52;
  assign rf_matrix_b_2_tile_v_3_MPORT_9_data = rf[rf_matrix_b_2_tile_v_3_MPORT_9_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_2_tile_v_2_MPORT_9_en = handshaked & _GEN_1393;
  assign rf_matrix_b_2_tile_v_2_MPORT_9_addr = 8'h56;
  assign rf_matrix_b_2_tile_v_2_MPORT_9_data = rf[rf_matrix_b_2_tile_v_2_MPORT_9_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_2_tile_v_1_MPORT_9_en = handshaked & _GEN_1393;
  assign rf_matrix_b_2_tile_v_1_MPORT_9_addr = 8'h5a;
  assign rf_matrix_b_2_tile_v_1_MPORT_9_data = rf[rf_matrix_b_2_tile_v_1_MPORT_9_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_2_tile_v_0_MPORT_9_en = handshaked & _GEN_1393;
  assign rf_matrix_b_2_tile_v_0_MPORT_9_addr = 8'h5e;
  assign rf_matrix_b_2_tile_v_0_MPORT_9_data = rf[rf_matrix_b_2_tile_v_0_MPORT_9_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_2_tile_v_3_MPORT_9_en = handshaked & _GEN_1393;
  assign rf_matrix_c_2_tile_v_3_MPORT_9_addr = 8'h83;
  assign rf_matrix_c_2_tile_v_3_MPORT_9_data = rf[rf_matrix_c_2_tile_v_3_MPORT_9_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_2_tile_v_2_MPORT_9_en = handshaked & _GEN_1393;
  assign rf_matrix_c_2_tile_v_2_MPORT_9_addr = 8'h87;
  assign rf_matrix_c_2_tile_v_2_MPORT_9_data = rf[rf_matrix_c_2_tile_v_2_MPORT_9_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_2_tile_v_1_MPORT_9_en = handshaked & _GEN_1393;
  assign rf_matrix_c_2_tile_v_1_MPORT_9_addr = 8'h8b;
  assign rf_matrix_c_2_tile_v_1_MPORT_9_data = rf[rf_matrix_c_2_tile_v_1_MPORT_9_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_2_tile_v_0_MPORT_9_en = handshaked & _GEN_1393;
  assign rf_matrix_c_2_tile_v_0_MPORT_9_addr = 8'h8f;
  assign rf_matrix_c_2_tile_v_0_MPORT_9_data = rf[rf_matrix_c_2_tile_v_0_MPORT_9_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_1_MPORT_58_en = handshaked & _GEN_1407;
  assign rf_a_tile_v_1_MPORT_58_addr = 8'h1;
  assign rf_a_tile_v_1_MPORT_58_data = rf[rf_a_tile_v_1_MPORT_58_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_0_MPORT_58_en = handshaked & _GEN_1407;
  assign rf_a_tile_v_0_MPORT_58_addr = 8'h5;
  assign rf_a_tile_v_0_MPORT_58_data = rf[rf_a_tile_v_0_MPORT_58_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_2_tile_v_3_MPORT_10_en = handshaked & _GEN_1407;
  assign rf_matrix_b_2_tile_v_3_MPORT_10_addr = 8'h52;
  assign rf_matrix_b_2_tile_v_3_MPORT_10_data = rf[rf_matrix_b_2_tile_v_3_MPORT_10_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_2_tile_v_2_MPORT_10_en = handshaked & _GEN_1407;
  assign rf_matrix_b_2_tile_v_2_MPORT_10_addr = 8'h56;
  assign rf_matrix_b_2_tile_v_2_MPORT_10_data = rf[rf_matrix_b_2_tile_v_2_MPORT_10_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_2_tile_v_1_MPORT_10_en = handshaked & _GEN_1407;
  assign rf_matrix_b_2_tile_v_1_MPORT_10_addr = 8'h5a;
  assign rf_matrix_b_2_tile_v_1_MPORT_10_data = rf[rf_matrix_b_2_tile_v_1_MPORT_10_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_2_tile_v_0_MPORT_10_en = handshaked & _GEN_1407;
  assign rf_matrix_b_2_tile_v_0_MPORT_10_addr = 8'h5e;
  assign rf_matrix_b_2_tile_v_0_MPORT_10_data = rf[rf_matrix_b_2_tile_v_0_MPORT_10_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_2_tile_v_3_MPORT_10_en = handshaked & _GEN_1407;
  assign rf_matrix_c_2_tile_v_3_MPORT_10_addr = 8'h86;
  assign rf_matrix_c_2_tile_v_3_MPORT_10_data = rf[rf_matrix_c_2_tile_v_3_MPORT_10_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_2_tile_v_2_MPORT_10_en = handshaked & _GEN_1407;
  assign rf_matrix_c_2_tile_v_2_MPORT_10_addr = 8'h87;
  assign rf_matrix_c_2_tile_v_2_MPORT_10_data = rf[rf_matrix_c_2_tile_v_2_MPORT_10_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_2_tile_v_1_MPORT_10_en = handshaked & _GEN_1407;
  assign rf_matrix_c_2_tile_v_1_MPORT_10_addr = 8'h8e;
  assign rf_matrix_c_2_tile_v_1_MPORT_10_data = rf[rf_matrix_c_2_tile_v_1_MPORT_10_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_2_tile_v_0_MPORT_10_en = handshaked & _GEN_1407;
  assign rf_matrix_c_2_tile_v_0_MPORT_10_addr = 8'h8f;
  assign rf_matrix_c_2_tile_v_0_MPORT_10_data = rf[rf_matrix_c_2_tile_v_0_MPORT_10_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_1_MPORT_59_en = handshaked & _GEN_1419;
  assign rf_a_tile_v_1_MPORT_59_addr = 8'h9;
  assign rf_a_tile_v_1_MPORT_59_data = rf[rf_a_tile_v_1_MPORT_59_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_0_MPORT_59_en = handshaked & _GEN_1419;
  assign rf_a_tile_v_0_MPORT_59_addr = 8'hd;
  assign rf_a_tile_v_0_MPORT_59_data = rf[rf_a_tile_v_0_MPORT_59_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_2_tile_v_3_MPORT_11_en = handshaked & _GEN_1419;
  assign rf_matrix_b_2_tile_v_3_MPORT_11_addr = 8'h52;
  assign rf_matrix_b_2_tile_v_3_MPORT_11_data = rf[rf_matrix_b_2_tile_v_3_MPORT_11_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_2_tile_v_2_MPORT_11_en = handshaked & _GEN_1419;
  assign rf_matrix_b_2_tile_v_2_MPORT_11_addr = 8'h56;
  assign rf_matrix_b_2_tile_v_2_MPORT_11_data = rf[rf_matrix_b_2_tile_v_2_MPORT_11_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_2_tile_v_1_MPORT_11_en = handshaked & _GEN_1419;
  assign rf_matrix_b_2_tile_v_1_MPORT_11_addr = 8'h5a;
  assign rf_matrix_b_2_tile_v_1_MPORT_11_data = rf[rf_matrix_b_2_tile_v_1_MPORT_11_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_2_tile_v_0_MPORT_11_en = handshaked & _GEN_1419;
  assign rf_matrix_b_2_tile_v_0_MPORT_11_addr = 8'h5e;
  assign rf_matrix_b_2_tile_v_0_MPORT_11_data = rf[rf_matrix_b_2_tile_v_0_MPORT_11_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_2_tile_v_3_MPORT_11_en = handshaked & _GEN_1419;
  assign rf_matrix_c_2_tile_v_3_MPORT_11_addr = 8'h96;
  assign rf_matrix_c_2_tile_v_3_MPORT_11_data = rf[rf_matrix_c_2_tile_v_3_MPORT_11_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_2_tile_v_2_MPORT_11_en = handshaked & _GEN_1419;
  assign rf_matrix_c_2_tile_v_2_MPORT_11_addr = 8'h97;
  assign rf_matrix_c_2_tile_v_2_MPORT_11_data = rf[rf_matrix_c_2_tile_v_2_MPORT_11_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_2_tile_v_1_MPORT_11_en = handshaked & _GEN_1419;
  assign rf_matrix_c_2_tile_v_1_MPORT_11_addr = 8'h9e;
  assign rf_matrix_c_2_tile_v_1_MPORT_11_data = rf[rf_matrix_c_2_tile_v_1_MPORT_11_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_2_tile_v_0_MPORT_11_en = handshaked & _GEN_1419;
  assign rf_matrix_c_2_tile_v_0_MPORT_11_addr = 8'h9f;
  assign rf_matrix_c_2_tile_v_0_MPORT_11_data = rf[rf_matrix_c_2_tile_v_0_MPORT_11_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_1_MPORT_60_en = handshaked & _GEN_1431;
  assign rf_a_tile_v_1_MPORT_60_addr = 8'h2;
  assign rf_a_tile_v_1_MPORT_60_data = rf[rf_a_tile_v_1_MPORT_60_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_0_MPORT_60_en = handshaked & _GEN_1431;
  assign rf_a_tile_v_0_MPORT_60_addr = 8'h6;
  assign rf_a_tile_v_0_MPORT_60_data = rf[rf_a_tile_v_0_MPORT_60_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_2_tile_v_3_MPORT_12_en = handshaked & _GEN_1431;
  assign rf_matrix_b_2_tile_v_3_MPORT_12_addr = 8'h62;
  assign rf_matrix_b_2_tile_v_3_MPORT_12_data = rf[rf_matrix_b_2_tile_v_3_MPORT_12_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_2_tile_v_2_MPORT_12_en = handshaked & _GEN_1431;
  assign rf_matrix_b_2_tile_v_2_MPORT_12_addr = 8'h66;
  assign rf_matrix_b_2_tile_v_2_MPORT_12_data = rf[rf_matrix_b_2_tile_v_2_MPORT_12_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_2_tile_v_1_MPORT_12_en = handshaked & _GEN_1431;
  assign rf_matrix_b_2_tile_v_1_MPORT_12_addr = 8'h6a;
  assign rf_matrix_b_2_tile_v_1_MPORT_12_data = rf[rf_matrix_b_2_tile_v_1_MPORT_12_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_2_tile_v_0_MPORT_12_en = handshaked & _GEN_1431;
  assign rf_matrix_b_2_tile_v_0_MPORT_12_addr = 8'h6e;
  assign rf_matrix_b_2_tile_v_0_MPORT_12_data = rf[rf_matrix_b_2_tile_v_0_MPORT_12_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_2_tile_v_3_MPORT_12_en = handshaked & _GEN_1431;
  assign rf_matrix_c_2_tile_v_3_MPORT_12_addr = 8'h84;
  assign rf_matrix_c_2_tile_v_3_MPORT_12_data = rf[rf_matrix_c_2_tile_v_3_MPORT_12_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_2_tile_v_2_MPORT_12_en = handshaked & _GEN_1431;
  assign rf_matrix_c_2_tile_v_2_MPORT_12_addr = 8'h85;
  assign rf_matrix_c_2_tile_v_2_MPORT_12_data = rf[rf_matrix_c_2_tile_v_2_MPORT_12_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_2_tile_v_1_MPORT_12_en = handshaked & _GEN_1431;
  assign rf_matrix_c_2_tile_v_1_MPORT_12_addr = 8'h8c;
  assign rf_matrix_c_2_tile_v_1_MPORT_12_data = rf[rf_matrix_c_2_tile_v_1_MPORT_12_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_2_tile_v_0_MPORT_12_en = handshaked & _GEN_1431;
  assign rf_matrix_c_2_tile_v_0_MPORT_12_addr = 8'h8d;
  assign rf_matrix_c_2_tile_v_0_MPORT_12_data = rf[rf_matrix_c_2_tile_v_0_MPORT_12_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_3_MPORT_20_en = handshaked & _GEN_1443;
  assign rf_a_tile_v_3_MPORT_20_addr = 8'h2;
  assign rf_a_tile_v_3_MPORT_20_data = rf[rf_a_tile_v_3_MPORT_20_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_2_MPORT_20_en = handshaked & _GEN_1443;
  assign rf_a_tile_v_2_MPORT_20_addr = 8'h6;
  assign rf_a_tile_v_2_MPORT_20_data = rf[rf_a_tile_v_2_MPORT_20_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_1_MPORT_61_en = handshaked & _GEN_1443;
  assign rf_a_tile_v_1_MPORT_61_addr = 8'ha;
  assign rf_a_tile_v_1_MPORT_61_data = rf[rf_a_tile_v_1_MPORT_61_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_0_MPORT_61_en = handshaked & _GEN_1443;
  assign rf_a_tile_v_0_MPORT_61_addr = 8'he;
  assign rf_a_tile_v_0_MPORT_61_data = rf[rf_a_tile_v_0_MPORT_61_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_2_tile_v_3_MPORT_13_en = handshaked & _GEN_1443;
  assign rf_matrix_b_2_tile_v_3_MPORT_13_addr = 8'h62;
  assign rf_matrix_b_2_tile_v_3_MPORT_13_data = rf[rf_matrix_b_2_tile_v_3_MPORT_13_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_2_tile_v_2_MPORT_13_en = handshaked & _GEN_1443;
  assign rf_matrix_b_2_tile_v_2_MPORT_13_addr = 8'h66;
  assign rf_matrix_b_2_tile_v_2_MPORT_13_data = rf[rf_matrix_b_2_tile_v_2_MPORT_13_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_2_tile_v_1_MPORT_13_en = handshaked & _GEN_1443;
  assign rf_matrix_b_2_tile_v_1_MPORT_13_addr = 8'h6a;
  assign rf_matrix_b_2_tile_v_1_MPORT_13_data = rf[rf_matrix_b_2_tile_v_1_MPORT_13_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_2_tile_v_0_MPORT_13_en = handshaked & _GEN_1443;
  assign rf_matrix_b_2_tile_v_0_MPORT_13_addr = 8'h6e;
  assign rf_matrix_b_2_tile_v_0_MPORT_13_data = rf[rf_matrix_b_2_tile_v_0_MPORT_13_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_2_tile_v_3_MPORT_13_en = handshaked & _GEN_1443;
  assign rf_matrix_c_2_tile_v_3_MPORT_13_addr = 8'h82;
  assign rf_matrix_c_2_tile_v_3_MPORT_13_data = rf[rf_matrix_c_2_tile_v_3_MPORT_13_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_2_tile_v_2_MPORT_13_en = handshaked & _GEN_1443;
  assign rf_matrix_c_2_tile_v_2_MPORT_13_addr = 8'h86;
  assign rf_matrix_c_2_tile_v_2_MPORT_13_data = rf[rf_matrix_c_2_tile_v_2_MPORT_13_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_2_tile_v_1_MPORT_13_en = handshaked & _GEN_1443;
  assign rf_matrix_c_2_tile_v_1_MPORT_13_addr = 8'h8a;
  assign rf_matrix_c_2_tile_v_1_MPORT_13_data = rf[rf_matrix_c_2_tile_v_1_MPORT_13_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_2_tile_v_0_MPORT_13_en = handshaked & _GEN_1443;
  assign rf_matrix_c_2_tile_v_0_MPORT_13_addr = 8'h8e;
  assign rf_matrix_c_2_tile_v_0_MPORT_13_data = rf[rf_matrix_c_2_tile_v_0_MPORT_13_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_1_MPORT_62_en = handshaked & _GEN_1457;
  assign rf_a_tile_v_1_MPORT_62_addr = 8'ha;
  assign rf_a_tile_v_1_MPORT_62_data = rf[rf_a_tile_v_1_MPORT_62_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_0_MPORT_62_en = handshaked & _GEN_1457;
  assign rf_a_tile_v_0_MPORT_62_addr = 8'he;
  assign rf_a_tile_v_0_MPORT_62_data = rf[rf_a_tile_v_0_MPORT_62_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_2_tile_v_3_MPORT_14_en = handshaked & _GEN_1457;
  assign rf_matrix_b_2_tile_v_3_MPORT_14_addr = 8'h62;
  assign rf_matrix_b_2_tile_v_3_MPORT_14_data = rf[rf_matrix_b_2_tile_v_3_MPORT_14_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_2_tile_v_2_MPORT_14_en = handshaked & _GEN_1457;
  assign rf_matrix_b_2_tile_v_2_MPORT_14_addr = 8'h66;
  assign rf_matrix_b_2_tile_v_2_MPORT_14_data = rf[rf_matrix_b_2_tile_v_2_MPORT_14_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_2_tile_v_1_MPORT_14_en = handshaked & _GEN_1457;
  assign rf_matrix_b_2_tile_v_1_MPORT_14_addr = 8'h6a;
  assign rf_matrix_b_2_tile_v_1_MPORT_14_data = rf[rf_matrix_b_2_tile_v_1_MPORT_14_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_2_tile_v_0_MPORT_14_en = handshaked & _GEN_1457;
  assign rf_matrix_b_2_tile_v_0_MPORT_14_addr = 8'h6e;
  assign rf_matrix_b_2_tile_v_0_MPORT_14_data = rf[rf_matrix_b_2_tile_v_0_MPORT_14_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_2_tile_v_3_MPORT_14_en = handshaked & _GEN_1457;
  assign rf_matrix_c_2_tile_v_3_MPORT_14_addr = 8'h94;
  assign rf_matrix_c_2_tile_v_3_MPORT_14_data = rf[rf_matrix_c_2_tile_v_3_MPORT_14_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_2_tile_v_2_MPORT_14_en = handshaked & _GEN_1457;
  assign rf_matrix_c_2_tile_v_2_MPORT_14_addr = 8'h95;
  assign rf_matrix_c_2_tile_v_2_MPORT_14_data = rf[rf_matrix_c_2_tile_v_2_MPORT_14_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_2_tile_v_1_MPORT_14_en = handshaked & _GEN_1457;
  assign rf_matrix_c_2_tile_v_1_MPORT_14_addr = 8'h9c;
  assign rf_matrix_c_2_tile_v_1_MPORT_14_data = rf[rf_matrix_c_2_tile_v_1_MPORT_14_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_2_tile_v_0_MPORT_14_en = handshaked & _GEN_1457;
  assign rf_matrix_c_2_tile_v_0_MPORT_14_addr = 8'h9d;
  assign rf_matrix_c_2_tile_v_0_MPORT_14_data = rf[rf_matrix_c_2_tile_v_0_MPORT_14_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_3_MPORT_21_en = handshaked & _GEN_1469;
  assign rf_a_tile_v_3_MPORT_21_addr = 8'h2;
  assign rf_a_tile_v_3_MPORT_21_data = rf[rf_a_tile_v_3_MPORT_21_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_2_MPORT_21_en = handshaked & _GEN_1469;
  assign rf_a_tile_v_2_MPORT_21_addr = 8'h6;
  assign rf_a_tile_v_2_MPORT_21_data = rf[rf_a_tile_v_2_MPORT_21_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_1_MPORT_63_en = handshaked & _GEN_1469;
  assign rf_a_tile_v_1_MPORT_63_addr = 8'ha;
  assign rf_a_tile_v_1_MPORT_63_data = rf[rf_a_tile_v_1_MPORT_63_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_0_MPORT_63_en = handshaked & _GEN_1469;
  assign rf_a_tile_v_0_MPORT_63_addr = 8'he;
  assign rf_a_tile_v_0_MPORT_63_data = rf[rf_a_tile_v_0_MPORT_63_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_2_tile_v_3_MPORT_15_en = handshaked & _GEN_1469;
  assign rf_matrix_b_2_tile_v_3_MPORT_15_addr = 8'h62;
  assign rf_matrix_b_2_tile_v_3_MPORT_15_data = rf[rf_matrix_b_2_tile_v_3_MPORT_15_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_2_tile_v_2_MPORT_15_en = handshaked & _GEN_1469;
  assign rf_matrix_b_2_tile_v_2_MPORT_15_addr = 8'h66;
  assign rf_matrix_b_2_tile_v_2_MPORT_15_data = rf[rf_matrix_b_2_tile_v_2_MPORT_15_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_2_tile_v_1_MPORT_15_en = handshaked & _GEN_1469;
  assign rf_matrix_b_2_tile_v_1_MPORT_15_addr = 8'h6a;
  assign rf_matrix_b_2_tile_v_1_MPORT_15_data = rf[rf_matrix_b_2_tile_v_1_MPORT_15_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_2_tile_v_0_MPORT_15_en = handshaked & _GEN_1469;
  assign rf_matrix_b_2_tile_v_0_MPORT_15_addr = 8'h6e;
  assign rf_matrix_b_2_tile_v_0_MPORT_15_data = rf[rf_matrix_b_2_tile_v_0_MPORT_15_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_2_tile_v_3_MPORT_15_en = handshaked & _GEN_1469;
  assign rf_matrix_c_2_tile_v_3_MPORT_15_addr = 8'h83;
  assign rf_matrix_c_2_tile_v_3_MPORT_15_data = rf[rf_matrix_c_2_tile_v_3_MPORT_15_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_2_tile_v_2_MPORT_15_en = handshaked & _GEN_1469;
  assign rf_matrix_c_2_tile_v_2_MPORT_15_addr = 8'h87;
  assign rf_matrix_c_2_tile_v_2_MPORT_15_data = rf[rf_matrix_c_2_tile_v_2_MPORT_15_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_2_tile_v_1_MPORT_15_en = handshaked & _GEN_1469;
  assign rf_matrix_c_2_tile_v_1_MPORT_15_addr = 8'h8b;
  assign rf_matrix_c_2_tile_v_1_MPORT_15_data = rf[rf_matrix_c_2_tile_v_1_MPORT_15_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_2_tile_v_0_MPORT_15_en = handshaked & _GEN_1469;
  assign rf_matrix_c_2_tile_v_0_MPORT_15_addr = 8'h8f;
  assign rf_matrix_c_2_tile_v_0_MPORT_15_data = rf[rf_matrix_c_2_tile_v_0_MPORT_15_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_1_MPORT_64_en = handshaked & _GEN_1483;
  assign rf_a_tile_v_1_MPORT_64_addr = 8'h2;
  assign rf_a_tile_v_1_MPORT_64_data = rf[rf_a_tile_v_1_MPORT_64_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_0_MPORT_64_en = handshaked & _GEN_1483;
  assign rf_a_tile_v_0_MPORT_64_addr = 8'h6;
  assign rf_a_tile_v_0_MPORT_64_data = rf[rf_a_tile_v_0_MPORT_64_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_2_tile_v_3_MPORT_16_en = handshaked & _GEN_1483;
  assign rf_matrix_b_2_tile_v_3_MPORT_16_addr = 8'h62;
  assign rf_matrix_b_2_tile_v_3_MPORT_16_data = rf[rf_matrix_b_2_tile_v_3_MPORT_16_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_2_tile_v_2_MPORT_16_en = handshaked & _GEN_1483;
  assign rf_matrix_b_2_tile_v_2_MPORT_16_addr = 8'h66;
  assign rf_matrix_b_2_tile_v_2_MPORT_16_data = rf[rf_matrix_b_2_tile_v_2_MPORT_16_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_2_tile_v_1_MPORT_16_en = handshaked & _GEN_1483;
  assign rf_matrix_b_2_tile_v_1_MPORT_16_addr = 8'h6a;
  assign rf_matrix_b_2_tile_v_1_MPORT_16_data = rf[rf_matrix_b_2_tile_v_1_MPORT_16_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_2_tile_v_0_MPORT_16_en = handshaked & _GEN_1483;
  assign rf_matrix_b_2_tile_v_0_MPORT_16_addr = 8'h6e;
  assign rf_matrix_b_2_tile_v_0_MPORT_16_data = rf[rf_matrix_b_2_tile_v_0_MPORT_16_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_2_tile_v_3_MPORT_16_en = handshaked & _GEN_1483;
  assign rf_matrix_c_2_tile_v_3_MPORT_16_addr = 8'h86;
  assign rf_matrix_c_2_tile_v_3_MPORT_16_data = rf[rf_matrix_c_2_tile_v_3_MPORT_16_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_2_tile_v_2_MPORT_16_en = handshaked & _GEN_1483;
  assign rf_matrix_c_2_tile_v_2_MPORT_16_addr = 8'h87;
  assign rf_matrix_c_2_tile_v_2_MPORT_16_data = rf[rf_matrix_c_2_tile_v_2_MPORT_16_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_2_tile_v_1_MPORT_16_en = handshaked & _GEN_1483;
  assign rf_matrix_c_2_tile_v_1_MPORT_16_addr = 8'h8e;
  assign rf_matrix_c_2_tile_v_1_MPORT_16_data = rf[rf_matrix_c_2_tile_v_1_MPORT_16_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_2_tile_v_0_MPORT_16_en = handshaked & _GEN_1483;
  assign rf_matrix_c_2_tile_v_0_MPORT_16_addr = 8'h8f;
  assign rf_matrix_c_2_tile_v_0_MPORT_16_data = rf[rf_matrix_c_2_tile_v_0_MPORT_16_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_1_MPORT_65_en = handshaked & _GEN_1495;
  assign rf_a_tile_v_1_MPORT_65_addr = 8'ha;
  assign rf_a_tile_v_1_MPORT_65_data = rf[rf_a_tile_v_1_MPORT_65_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_0_MPORT_65_en = handshaked & _GEN_1495;
  assign rf_a_tile_v_0_MPORT_65_addr = 8'he;
  assign rf_a_tile_v_0_MPORT_65_data = rf[rf_a_tile_v_0_MPORT_65_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_2_tile_v_3_MPORT_17_en = handshaked & _GEN_1495;
  assign rf_matrix_b_2_tile_v_3_MPORT_17_addr = 8'h62;
  assign rf_matrix_b_2_tile_v_3_MPORT_17_data = rf[rf_matrix_b_2_tile_v_3_MPORT_17_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_2_tile_v_2_MPORT_17_en = handshaked & _GEN_1495;
  assign rf_matrix_b_2_tile_v_2_MPORT_17_addr = 8'h66;
  assign rf_matrix_b_2_tile_v_2_MPORT_17_data = rf[rf_matrix_b_2_tile_v_2_MPORT_17_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_2_tile_v_1_MPORT_17_en = handshaked & _GEN_1495;
  assign rf_matrix_b_2_tile_v_1_MPORT_17_addr = 8'h6a;
  assign rf_matrix_b_2_tile_v_1_MPORT_17_data = rf[rf_matrix_b_2_tile_v_1_MPORT_17_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_2_tile_v_0_MPORT_17_en = handshaked & _GEN_1495;
  assign rf_matrix_b_2_tile_v_0_MPORT_17_addr = 8'h6e;
  assign rf_matrix_b_2_tile_v_0_MPORT_17_data = rf[rf_matrix_b_2_tile_v_0_MPORT_17_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_2_tile_v_3_MPORT_17_en = handshaked & _GEN_1495;
  assign rf_matrix_c_2_tile_v_3_MPORT_17_addr = 8'h96;
  assign rf_matrix_c_2_tile_v_3_MPORT_17_data = rf[rf_matrix_c_2_tile_v_3_MPORT_17_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_2_tile_v_2_MPORT_17_en = handshaked & _GEN_1495;
  assign rf_matrix_c_2_tile_v_2_MPORT_17_addr = 8'h97;
  assign rf_matrix_c_2_tile_v_2_MPORT_17_data = rf[rf_matrix_c_2_tile_v_2_MPORT_17_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_2_tile_v_1_MPORT_17_en = handshaked & _GEN_1495;
  assign rf_matrix_c_2_tile_v_1_MPORT_17_addr = 8'h9e;
  assign rf_matrix_c_2_tile_v_1_MPORT_17_data = rf[rf_matrix_c_2_tile_v_1_MPORT_17_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_2_tile_v_0_MPORT_17_en = handshaked & _GEN_1495;
  assign rf_matrix_c_2_tile_v_0_MPORT_17_addr = 8'h9f;
  assign rf_matrix_c_2_tile_v_0_MPORT_17_data = rf[rf_matrix_c_2_tile_v_0_MPORT_17_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_1_MPORT_66_en = handshaked & _GEN_1507;
  assign rf_a_tile_v_1_MPORT_66_addr = 8'h3;
  assign rf_a_tile_v_1_MPORT_66_data = rf[rf_a_tile_v_1_MPORT_66_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_0_MPORT_66_en = handshaked & _GEN_1507;
  assign rf_a_tile_v_0_MPORT_66_addr = 8'h7;
  assign rf_a_tile_v_0_MPORT_66_data = rf[rf_a_tile_v_0_MPORT_66_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_2_tile_v_3_MPORT_18_en = handshaked & _GEN_1507;
  assign rf_matrix_b_2_tile_v_3_MPORT_18_addr = 8'h72;
  assign rf_matrix_b_2_tile_v_3_MPORT_18_data = rf[rf_matrix_b_2_tile_v_3_MPORT_18_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_2_tile_v_2_MPORT_18_en = handshaked & _GEN_1507;
  assign rf_matrix_b_2_tile_v_2_MPORT_18_addr = 8'h76;
  assign rf_matrix_b_2_tile_v_2_MPORT_18_data = rf[rf_matrix_b_2_tile_v_2_MPORT_18_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_2_tile_v_1_MPORT_18_en = handshaked & _GEN_1507;
  assign rf_matrix_b_2_tile_v_1_MPORT_18_addr = 8'h7a;
  assign rf_matrix_b_2_tile_v_1_MPORT_18_data = rf[rf_matrix_b_2_tile_v_1_MPORT_18_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_2_tile_v_0_MPORT_18_en = handshaked & _GEN_1507;
  assign rf_matrix_b_2_tile_v_0_MPORT_18_addr = 8'h7e;
  assign rf_matrix_b_2_tile_v_0_MPORT_18_data = rf[rf_matrix_b_2_tile_v_0_MPORT_18_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_2_tile_v_3_MPORT_18_en = handshaked & _GEN_1507;
  assign rf_matrix_c_2_tile_v_3_MPORT_18_addr = 8'h84;
  assign rf_matrix_c_2_tile_v_3_MPORT_18_data = rf[rf_matrix_c_2_tile_v_3_MPORT_18_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_2_tile_v_2_MPORT_18_en = handshaked & _GEN_1507;
  assign rf_matrix_c_2_tile_v_2_MPORT_18_addr = 8'h85;
  assign rf_matrix_c_2_tile_v_2_MPORT_18_data = rf[rf_matrix_c_2_tile_v_2_MPORT_18_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_2_tile_v_1_MPORT_18_en = handshaked & _GEN_1507;
  assign rf_matrix_c_2_tile_v_1_MPORT_18_addr = 8'h8c;
  assign rf_matrix_c_2_tile_v_1_MPORT_18_data = rf[rf_matrix_c_2_tile_v_1_MPORT_18_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_2_tile_v_0_MPORT_18_en = handshaked & _GEN_1507;
  assign rf_matrix_c_2_tile_v_0_MPORT_18_addr = 8'h8d;
  assign rf_matrix_c_2_tile_v_0_MPORT_18_data = rf[rf_matrix_c_2_tile_v_0_MPORT_18_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_3_MPORT_22_en = handshaked & _GEN_1519;
  assign rf_a_tile_v_3_MPORT_22_addr = 8'h3;
  assign rf_a_tile_v_3_MPORT_22_data = rf[rf_a_tile_v_3_MPORT_22_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_2_MPORT_22_en = handshaked & _GEN_1519;
  assign rf_a_tile_v_2_MPORT_22_addr = 8'h7;
  assign rf_a_tile_v_2_MPORT_22_data = rf[rf_a_tile_v_2_MPORT_22_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_1_MPORT_67_en = handshaked & _GEN_1519;
  assign rf_a_tile_v_1_MPORT_67_addr = 8'hb;
  assign rf_a_tile_v_1_MPORT_67_data = rf[rf_a_tile_v_1_MPORT_67_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_0_MPORT_67_en = handshaked & _GEN_1519;
  assign rf_a_tile_v_0_MPORT_67_addr = 8'hf;
  assign rf_a_tile_v_0_MPORT_67_data = rf[rf_a_tile_v_0_MPORT_67_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_2_tile_v_3_MPORT_19_en = handshaked & _GEN_1519;
  assign rf_matrix_b_2_tile_v_3_MPORT_19_addr = 8'h72;
  assign rf_matrix_b_2_tile_v_3_MPORT_19_data = rf[rf_matrix_b_2_tile_v_3_MPORT_19_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_2_tile_v_2_MPORT_19_en = handshaked & _GEN_1519;
  assign rf_matrix_b_2_tile_v_2_MPORT_19_addr = 8'h76;
  assign rf_matrix_b_2_tile_v_2_MPORT_19_data = rf[rf_matrix_b_2_tile_v_2_MPORT_19_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_2_tile_v_1_MPORT_19_en = handshaked & _GEN_1519;
  assign rf_matrix_b_2_tile_v_1_MPORT_19_addr = 8'h7a;
  assign rf_matrix_b_2_tile_v_1_MPORT_19_data = rf[rf_matrix_b_2_tile_v_1_MPORT_19_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_2_tile_v_0_MPORT_19_en = handshaked & _GEN_1519;
  assign rf_matrix_b_2_tile_v_0_MPORT_19_addr = 8'h7e;
  assign rf_matrix_b_2_tile_v_0_MPORT_19_data = rf[rf_matrix_b_2_tile_v_0_MPORT_19_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_2_tile_v_3_MPORT_19_en = handshaked & _GEN_1519;
  assign rf_matrix_c_2_tile_v_3_MPORT_19_addr = 8'h82;
  assign rf_matrix_c_2_tile_v_3_MPORT_19_data = rf[rf_matrix_c_2_tile_v_3_MPORT_19_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_2_tile_v_2_MPORT_19_en = handshaked & _GEN_1519;
  assign rf_matrix_c_2_tile_v_2_MPORT_19_addr = 8'h86;
  assign rf_matrix_c_2_tile_v_2_MPORT_19_data = rf[rf_matrix_c_2_tile_v_2_MPORT_19_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_2_tile_v_1_MPORT_19_en = handshaked & _GEN_1519;
  assign rf_matrix_c_2_tile_v_1_MPORT_19_addr = 8'h8a;
  assign rf_matrix_c_2_tile_v_1_MPORT_19_data = rf[rf_matrix_c_2_tile_v_1_MPORT_19_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_2_tile_v_0_MPORT_19_en = handshaked & _GEN_1519;
  assign rf_matrix_c_2_tile_v_0_MPORT_19_addr = 8'h8e;
  assign rf_matrix_c_2_tile_v_0_MPORT_19_data = rf[rf_matrix_c_2_tile_v_0_MPORT_19_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_1_MPORT_68_en = handshaked & _GEN_1533;
  assign rf_a_tile_v_1_MPORT_68_addr = 8'hb;
  assign rf_a_tile_v_1_MPORT_68_data = rf[rf_a_tile_v_1_MPORT_68_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_0_MPORT_68_en = handshaked & _GEN_1533;
  assign rf_a_tile_v_0_MPORT_68_addr = 8'hf;
  assign rf_a_tile_v_0_MPORT_68_data = rf[rf_a_tile_v_0_MPORT_68_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_2_tile_v_3_MPORT_20_en = handshaked & _GEN_1533;
  assign rf_matrix_b_2_tile_v_3_MPORT_20_addr = 8'h72;
  assign rf_matrix_b_2_tile_v_3_MPORT_20_data = rf[rf_matrix_b_2_tile_v_3_MPORT_20_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_2_tile_v_2_MPORT_20_en = handshaked & _GEN_1533;
  assign rf_matrix_b_2_tile_v_2_MPORT_20_addr = 8'h76;
  assign rf_matrix_b_2_tile_v_2_MPORT_20_data = rf[rf_matrix_b_2_tile_v_2_MPORT_20_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_2_tile_v_1_MPORT_20_en = handshaked & _GEN_1533;
  assign rf_matrix_b_2_tile_v_1_MPORT_20_addr = 8'h7a;
  assign rf_matrix_b_2_tile_v_1_MPORT_20_data = rf[rf_matrix_b_2_tile_v_1_MPORT_20_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_2_tile_v_0_MPORT_20_en = handshaked & _GEN_1533;
  assign rf_matrix_b_2_tile_v_0_MPORT_20_addr = 8'h7e;
  assign rf_matrix_b_2_tile_v_0_MPORT_20_data = rf[rf_matrix_b_2_tile_v_0_MPORT_20_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_2_tile_v_3_MPORT_20_en = handshaked & _GEN_1533;
  assign rf_matrix_c_2_tile_v_3_MPORT_20_addr = 8'h94;
  assign rf_matrix_c_2_tile_v_3_MPORT_20_data = rf[rf_matrix_c_2_tile_v_3_MPORT_20_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_2_tile_v_2_MPORT_20_en = handshaked & _GEN_1533;
  assign rf_matrix_c_2_tile_v_2_MPORT_20_addr = 8'h95;
  assign rf_matrix_c_2_tile_v_2_MPORT_20_data = rf[rf_matrix_c_2_tile_v_2_MPORT_20_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_2_tile_v_1_MPORT_20_en = handshaked & _GEN_1533;
  assign rf_matrix_c_2_tile_v_1_MPORT_20_addr = 8'h9c;
  assign rf_matrix_c_2_tile_v_1_MPORT_20_data = rf[rf_matrix_c_2_tile_v_1_MPORT_20_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_2_tile_v_0_MPORT_20_en = handshaked & _GEN_1533;
  assign rf_matrix_c_2_tile_v_0_MPORT_20_addr = 8'h9d;
  assign rf_matrix_c_2_tile_v_0_MPORT_20_data = rf[rf_matrix_c_2_tile_v_0_MPORT_20_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_3_MPORT_23_en = handshaked & _GEN_1545;
  assign rf_a_tile_v_3_MPORT_23_addr = 8'h3;
  assign rf_a_tile_v_3_MPORT_23_data = rf[rf_a_tile_v_3_MPORT_23_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_2_MPORT_23_en = handshaked & _GEN_1545;
  assign rf_a_tile_v_2_MPORT_23_addr = 8'h7;
  assign rf_a_tile_v_2_MPORT_23_data = rf[rf_a_tile_v_2_MPORT_23_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_1_MPORT_69_en = handshaked & _GEN_1545;
  assign rf_a_tile_v_1_MPORT_69_addr = 8'hb;
  assign rf_a_tile_v_1_MPORT_69_data = rf[rf_a_tile_v_1_MPORT_69_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_0_MPORT_69_en = handshaked & _GEN_1545;
  assign rf_a_tile_v_0_MPORT_69_addr = 8'hf;
  assign rf_a_tile_v_0_MPORT_69_data = rf[rf_a_tile_v_0_MPORT_69_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_2_tile_v_3_MPORT_21_en = handshaked & _GEN_1545;
  assign rf_matrix_b_2_tile_v_3_MPORT_21_addr = 8'h72;
  assign rf_matrix_b_2_tile_v_3_MPORT_21_data = rf[rf_matrix_b_2_tile_v_3_MPORT_21_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_2_tile_v_2_MPORT_21_en = handshaked & _GEN_1545;
  assign rf_matrix_b_2_tile_v_2_MPORT_21_addr = 8'h76;
  assign rf_matrix_b_2_tile_v_2_MPORT_21_data = rf[rf_matrix_b_2_tile_v_2_MPORT_21_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_2_tile_v_1_MPORT_21_en = handshaked & _GEN_1545;
  assign rf_matrix_b_2_tile_v_1_MPORT_21_addr = 8'h7a;
  assign rf_matrix_b_2_tile_v_1_MPORT_21_data = rf[rf_matrix_b_2_tile_v_1_MPORT_21_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_2_tile_v_0_MPORT_21_en = handshaked & _GEN_1545;
  assign rf_matrix_b_2_tile_v_0_MPORT_21_addr = 8'h7e;
  assign rf_matrix_b_2_tile_v_0_MPORT_21_data = rf[rf_matrix_b_2_tile_v_0_MPORT_21_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_2_tile_v_3_MPORT_21_en = handshaked & _GEN_1545;
  assign rf_matrix_c_2_tile_v_3_MPORT_21_addr = 8'h83;
  assign rf_matrix_c_2_tile_v_3_MPORT_21_data = rf[rf_matrix_c_2_tile_v_3_MPORT_21_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_2_tile_v_2_MPORT_21_en = handshaked & _GEN_1545;
  assign rf_matrix_c_2_tile_v_2_MPORT_21_addr = 8'h87;
  assign rf_matrix_c_2_tile_v_2_MPORT_21_data = rf[rf_matrix_c_2_tile_v_2_MPORT_21_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_2_tile_v_1_MPORT_21_en = handshaked & _GEN_1545;
  assign rf_matrix_c_2_tile_v_1_MPORT_21_addr = 8'h8b;
  assign rf_matrix_c_2_tile_v_1_MPORT_21_data = rf[rf_matrix_c_2_tile_v_1_MPORT_21_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_2_tile_v_0_MPORT_21_en = handshaked & _GEN_1545;
  assign rf_matrix_c_2_tile_v_0_MPORT_21_addr = 8'h8f;
  assign rf_matrix_c_2_tile_v_0_MPORT_21_data = rf[rf_matrix_c_2_tile_v_0_MPORT_21_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_1_MPORT_70_en = handshaked & _GEN_1559;
  assign rf_a_tile_v_1_MPORT_70_addr = 8'h3;
  assign rf_a_tile_v_1_MPORT_70_data = rf[rf_a_tile_v_1_MPORT_70_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_0_MPORT_70_en = handshaked & _GEN_1559;
  assign rf_a_tile_v_0_MPORT_70_addr = 8'h7;
  assign rf_a_tile_v_0_MPORT_70_data = rf[rf_a_tile_v_0_MPORT_70_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_2_tile_v_3_MPORT_22_en = handshaked & _GEN_1559;
  assign rf_matrix_b_2_tile_v_3_MPORT_22_addr = 8'h72;
  assign rf_matrix_b_2_tile_v_3_MPORT_22_data = rf[rf_matrix_b_2_tile_v_3_MPORT_22_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_2_tile_v_2_MPORT_22_en = handshaked & _GEN_1559;
  assign rf_matrix_b_2_tile_v_2_MPORT_22_addr = 8'h76;
  assign rf_matrix_b_2_tile_v_2_MPORT_22_data = rf[rf_matrix_b_2_tile_v_2_MPORT_22_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_2_tile_v_1_MPORT_22_en = handshaked & _GEN_1559;
  assign rf_matrix_b_2_tile_v_1_MPORT_22_addr = 8'h7a;
  assign rf_matrix_b_2_tile_v_1_MPORT_22_data = rf[rf_matrix_b_2_tile_v_1_MPORT_22_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_2_tile_v_0_MPORT_22_en = handshaked & _GEN_1559;
  assign rf_matrix_b_2_tile_v_0_MPORT_22_addr = 8'h7e;
  assign rf_matrix_b_2_tile_v_0_MPORT_22_data = rf[rf_matrix_b_2_tile_v_0_MPORT_22_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_2_tile_v_3_MPORT_22_en = handshaked & _GEN_1559;
  assign rf_matrix_c_2_tile_v_3_MPORT_22_addr = 8'h86;
  assign rf_matrix_c_2_tile_v_3_MPORT_22_data = rf[rf_matrix_c_2_tile_v_3_MPORT_22_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_2_tile_v_2_MPORT_22_en = handshaked & _GEN_1559;
  assign rf_matrix_c_2_tile_v_2_MPORT_22_addr = 8'h87;
  assign rf_matrix_c_2_tile_v_2_MPORT_22_data = rf[rf_matrix_c_2_tile_v_2_MPORT_22_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_2_tile_v_1_MPORT_22_en = handshaked & _GEN_1559;
  assign rf_matrix_c_2_tile_v_1_MPORT_22_addr = 8'h8e;
  assign rf_matrix_c_2_tile_v_1_MPORT_22_data = rf[rf_matrix_c_2_tile_v_1_MPORT_22_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_2_tile_v_0_MPORT_22_en = handshaked & _GEN_1559;
  assign rf_matrix_c_2_tile_v_0_MPORT_22_addr = 8'h8f;
  assign rf_matrix_c_2_tile_v_0_MPORT_22_data = rf[rf_matrix_c_2_tile_v_0_MPORT_22_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_1_MPORT_71_en = handshaked & _GEN_1571;
  assign rf_a_tile_v_1_MPORT_71_addr = 8'hb;
  assign rf_a_tile_v_1_MPORT_71_data = rf[rf_a_tile_v_1_MPORT_71_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_0_MPORT_71_en = handshaked & _GEN_1571;
  assign rf_a_tile_v_0_MPORT_71_addr = 8'hf;
  assign rf_a_tile_v_0_MPORT_71_data = rf[rf_a_tile_v_0_MPORT_71_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_2_tile_v_3_MPORT_23_en = handshaked & _GEN_1571;
  assign rf_matrix_b_2_tile_v_3_MPORT_23_addr = 8'h72;
  assign rf_matrix_b_2_tile_v_3_MPORT_23_data = rf[rf_matrix_b_2_tile_v_3_MPORT_23_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_2_tile_v_2_MPORT_23_en = handshaked & _GEN_1571;
  assign rf_matrix_b_2_tile_v_2_MPORT_23_addr = 8'h76;
  assign rf_matrix_b_2_tile_v_2_MPORT_23_data = rf[rf_matrix_b_2_tile_v_2_MPORT_23_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_2_tile_v_1_MPORT_23_en = handshaked & _GEN_1571;
  assign rf_matrix_b_2_tile_v_1_MPORT_23_addr = 8'h7a;
  assign rf_matrix_b_2_tile_v_1_MPORT_23_data = rf[rf_matrix_b_2_tile_v_1_MPORT_23_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_2_tile_v_0_MPORT_23_en = handshaked & _GEN_1571;
  assign rf_matrix_b_2_tile_v_0_MPORT_23_addr = 8'h7e;
  assign rf_matrix_b_2_tile_v_0_MPORT_23_data = rf[rf_matrix_b_2_tile_v_0_MPORT_23_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_2_tile_v_3_MPORT_23_en = handshaked & _GEN_1571;
  assign rf_matrix_c_2_tile_v_3_MPORT_23_addr = 8'h96;
  assign rf_matrix_c_2_tile_v_3_MPORT_23_data = rf[rf_matrix_c_2_tile_v_3_MPORT_23_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_2_tile_v_2_MPORT_23_en = handshaked & _GEN_1571;
  assign rf_matrix_c_2_tile_v_2_MPORT_23_addr = 8'h97;
  assign rf_matrix_c_2_tile_v_2_MPORT_23_data = rf[rf_matrix_c_2_tile_v_2_MPORT_23_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_2_tile_v_1_MPORT_23_en = handshaked & _GEN_1571;
  assign rf_matrix_c_2_tile_v_1_MPORT_23_addr = 8'h9e;
  assign rf_matrix_c_2_tile_v_1_MPORT_23_data = rf[rf_matrix_c_2_tile_v_1_MPORT_23_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_2_tile_v_0_MPORT_23_en = handshaked & _GEN_1571;
  assign rf_matrix_c_2_tile_v_0_MPORT_23_addr = 8'h9f;
  assign rf_matrix_c_2_tile_v_0_MPORT_23_data = rf[rf_matrix_c_2_tile_v_0_MPORT_23_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_1_MPORT_72_en = handshaked & _GEN_1276;
  assign rf_a_tile_v_1_MPORT_72_addr = 8'h20;
  assign rf_a_tile_v_1_MPORT_72_data = rf[rf_a_tile_v_1_MPORT_72_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_0_MPORT_72_en = handshaked & _GEN_1276;
  assign rf_a_tile_v_0_MPORT_72_addr = 8'h24;
  assign rf_a_tile_v_0_MPORT_72_data = rf[rf_a_tile_v_0_MPORT_72_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_3_tile_v_3_MPORT_en = handshaked & _GEN_1276;
  assign rf_matrix_b_3_tile_v_3_MPORT_addr = 8'h42;
  assign rf_matrix_b_3_tile_v_3_MPORT_data = rf[rf_matrix_b_3_tile_v_3_MPORT_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_3_tile_v_2_MPORT_en = handshaked & _GEN_1276;
  assign rf_matrix_b_3_tile_v_2_MPORT_addr = 8'h46;
  assign rf_matrix_b_3_tile_v_2_MPORT_data = rf[rf_matrix_b_3_tile_v_2_MPORT_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_3_tile_v_1_MPORT_en = handshaked & _GEN_1276;
  assign rf_matrix_b_3_tile_v_1_MPORT_addr = 8'h4a;
  assign rf_matrix_b_3_tile_v_1_MPORT_data = rf[rf_matrix_b_3_tile_v_1_MPORT_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_3_tile_v_0_MPORT_en = handshaked & _GEN_1276;
  assign rf_matrix_b_3_tile_v_0_MPORT_addr = 8'h4e;
  assign rf_matrix_b_3_tile_v_0_MPORT_data = rf[rf_matrix_b_3_tile_v_0_MPORT_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_3_tile_v_3_MPORT_en = handshaked & _GEN_1276;
  assign rf_matrix_c_3_tile_v_3_MPORT_addr = 8'hc4;
  assign rf_matrix_c_3_tile_v_3_MPORT_data = rf[rf_matrix_c_3_tile_v_3_MPORT_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_3_tile_v_2_MPORT_en = handshaked & _GEN_1276;
  assign rf_matrix_c_3_tile_v_2_MPORT_addr = 8'hc5;
  assign rf_matrix_c_3_tile_v_2_MPORT_data = rf[rf_matrix_c_3_tile_v_2_MPORT_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_3_tile_v_1_MPORT_en = handshaked & _GEN_1276;
  assign rf_matrix_c_3_tile_v_1_MPORT_addr = 8'hcc;
  assign rf_matrix_c_3_tile_v_1_MPORT_data = rf[rf_matrix_c_3_tile_v_1_MPORT_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_3_tile_v_0_MPORT_en = handshaked & _GEN_1276;
  assign rf_matrix_c_3_tile_v_0_MPORT_addr = 8'hcd;
  assign rf_matrix_c_3_tile_v_0_MPORT_data = rf[rf_matrix_c_3_tile_v_0_MPORT_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_3_MPORT_24_en = handshaked & _GEN_1291;
  assign rf_a_tile_v_3_MPORT_24_addr = 8'h20;
  assign rf_a_tile_v_3_MPORT_24_data = rf[rf_a_tile_v_3_MPORT_24_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_2_MPORT_24_en = handshaked & _GEN_1291;
  assign rf_a_tile_v_2_MPORT_24_addr = 8'h24;
  assign rf_a_tile_v_2_MPORT_24_data = rf[rf_a_tile_v_2_MPORT_24_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_1_MPORT_73_en = handshaked & _GEN_1291;
  assign rf_a_tile_v_1_MPORT_73_addr = 8'h28;
  assign rf_a_tile_v_1_MPORT_73_data = rf[rf_a_tile_v_1_MPORT_73_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_0_MPORT_73_en = handshaked & _GEN_1291;
  assign rf_a_tile_v_0_MPORT_73_addr = 8'h2c;
  assign rf_a_tile_v_0_MPORT_73_data = rf[rf_a_tile_v_0_MPORT_73_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_3_tile_v_3_MPORT_1_en = handshaked & _GEN_1291;
  assign rf_matrix_b_3_tile_v_3_MPORT_1_addr = 8'h42;
  assign rf_matrix_b_3_tile_v_3_MPORT_1_data = rf[rf_matrix_b_3_tile_v_3_MPORT_1_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_3_tile_v_2_MPORT_1_en = handshaked & _GEN_1291;
  assign rf_matrix_b_3_tile_v_2_MPORT_1_addr = 8'h46;
  assign rf_matrix_b_3_tile_v_2_MPORT_1_data = rf[rf_matrix_b_3_tile_v_2_MPORT_1_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_3_tile_v_1_MPORT_1_en = handshaked & _GEN_1291;
  assign rf_matrix_b_3_tile_v_1_MPORT_1_addr = 8'h4a;
  assign rf_matrix_b_3_tile_v_1_MPORT_1_data = rf[rf_matrix_b_3_tile_v_1_MPORT_1_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_3_tile_v_0_MPORT_1_en = handshaked & _GEN_1291;
  assign rf_matrix_b_3_tile_v_0_MPORT_1_addr = 8'h4e;
  assign rf_matrix_b_3_tile_v_0_MPORT_1_data = rf[rf_matrix_b_3_tile_v_0_MPORT_1_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_3_tile_v_3_MPORT_1_en = handshaked & _GEN_1291;
  assign rf_matrix_c_3_tile_v_3_MPORT_1_addr = 8'ha2;
  assign rf_matrix_c_3_tile_v_3_MPORT_1_data = rf[rf_matrix_c_3_tile_v_3_MPORT_1_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_3_tile_v_2_MPORT_1_en = handshaked & _GEN_1291;
  assign rf_matrix_c_3_tile_v_2_MPORT_1_addr = 8'ha6;
  assign rf_matrix_c_3_tile_v_2_MPORT_1_data = rf[rf_matrix_c_3_tile_v_2_MPORT_1_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_3_tile_v_1_MPORT_1_en = handshaked & _GEN_1291;
  assign rf_matrix_c_3_tile_v_1_MPORT_1_addr = 8'haa;
  assign rf_matrix_c_3_tile_v_1_MPORT_1_data = rf[rf_matrix_c_3_tile_v_1_MPORT_1_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_3_tile_v_0_MPORT_1_en = handshaked & _GEN_1291;
  assign rf_matrix_c_3_tile_v_0_MPORT_1_addr = 8'hae;
  assign rf_matrix_c_3_tile_v_0_MPORT_1_data = rf[rf_matrix_c_3_tile_v_0_MPORT_1_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_1_MPORT_74_en = handshaked & _GEN_1305;
  assign rf_a_tile_v_1_MPORT_74_addr = 8'h28;
  assign rf_a_tile_v_1_MPORT_74_data = rf[rf_a_tile_v_1_MPORT_74_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_0_MPORT_74_en = handshaked & _GEN_1305;
  assign rf_a_tile_v_0_MPORT_74_addr = 8'h2c;
  assign rf_a_tile_v_0_MPORT_74_data = rf[rf_a_tile_v_0_MPORT_74_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_3_tile_v_3_MPORT_2_en = handshaked & _GEN_1305;
  assign rf_matrix_b_3_tile_v_3_MPORT_2_addr = 8'h42;
  assign rf_matrix_b_3_tile_v_3_MPORT_2_data = rf[rf_matrix_b_3_tile_v_3_MPORT_2_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_3_tile_v_2_MPORT_2_en = handshaked & _GEN_1305;
  assign rf_matrix_b_3_tile_v_2_MPORT_2_addr = 8'h46;
  assign rf_matrix_b_3_tile_v_2_MPORT_2_data = rf[rf_matrix_b_3_tile_v_2_MPORT_2_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_3_tile_v_1_MPORT_2_en = handshaked & _GEN_1305;
  assign rf_matrix_b_3_tile_v_1_MPORT_2_addr = 8'h4a;
  assign rf_matrix_b_3_tile_v_1_MPORT_2_data = rf[rf_matrix_b_3_tile_v_1_MPORT_2_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_3_tile_v_0_MPORT_2_en = handshaked & _GEN_1305;
  assign rf_matrix_b_3_tile_v_0_MPORT_2_addr = 8'h4e;
  assign rf_matrix_b_3_tile_v_0_MPORT_2_data = rf[rf_matrix_b_3_tile_v_0_MPORT_2_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_3_tile_v_3_MPORT_2_en = handshaked & _GEN_1305;
  assign rf_matrix_c_3_tile_v_3_MPORT_2_addr = 8'hd4;
  assign rf_matrix_c_3_tile_v_3_MPORT_2_data = rf[rf_matrix_c_3_tile_v_3_MPORT_2_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_3_tile_v_2_MPORT_2_en = handshaked & _GEN_1305;
  assign rf_matrix_c_3_tile_v_2_MPORT_2_addr = 8'hd5;
  assign rf_matrix_c_3_tile_v_2_MPORT_2_data = rf[rf_matrix_c_3_tile_v_2_MPORT_2_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_3_tile_v_1_MPORT_2_en = handshaked & _GEN_1305;
  assign rf_matrix_c_3_tile_v_1_MPORT_2_addr = 8'hdc;
  assign rf_matrix_c_3_tile_v_1_MPORT_2_data = rf[rf_matrix_c_3_tile_v_1_MPORT_2_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_3_tile_v_0_MPORT_2_en = handshaked & _GEN_1305;
  assign rf_matrix_c_3_tile_v_0_MPORT_2_addr = 8'hdd;
  assign rf_matrix_c_3_tile_v_0_MPORT_2_data = rf[rf_matrix_c_3_tile_v_0_MPORT_2_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_3_MPORT_25_en = handshaked & _GEN_1317;
  assign rf_a_tile_v_3_MPORT_25_addr = 8'h20;
  assign rf_a_tile_v_3_MPORT_25_data = rf[rf_a_tile_v_3_MPORT_25_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_2_MPORT_25_en = handshaked & _GEN_1317;
  assign rf_a_tile_v_2_MPORT_25_addr = 8'h24;
  assign rf_a_tile_v_2_MPORT_25_data = rf[rf_a_tile_v_2_MPORT_25_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_1_MPORT_75_en = handshaked & _GEN_1317;
  assign rf_a_tile_v_1_MPORT_75_addr = 8'h28;
  assign rf_a_tile_v_1_MPORT_75_data = rf[rf_a_tile_v_1_MPORT_75_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_0_MPORT_75_en = handshaked & _GEN_1317;
  assign rf_a_tile_v_0_MPORT_75_addr = 8'h2c;
  assign rf_a_tile_v_0_MPORT_75_data = rf[rf_a_tile_v_0_MPORT_75_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_3_tile_v_3_MPORT_3_en = handshaked & _GEN_1317;
  assign rf_matrix_b_3_tile_v_3_MPORT_3_addr = 8'h42;
  assign rf_matrix_b_3_tile_v_3_MPORT_3_data = rf[rf_matrix_b_3_tile_v_3_MPORT_3_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_3_tile_v_2_MPORT_3_en = handshaked & _GEN_1317;
  assign rf_matrix_b_3_tile_v_2_MPORT_3_addr = 8'h46;
  assign rf_matrix_b_3_tile_v_2_MPORT_3_data = rf[rf_matrix_b_3_tile_v_2_MPORT_3_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_3_tile_v_1_MPORT_3_en = handshaked & _GEN_1317;
  assign rf_matrix_b_3_tile_v_1_MPORT_3_addr = 8'h4a;
  assign rf_matrix_b_3_tile_v_1_MPORT_3_data = rf[rf_matrix_b_3_tile_v_1_MPORT_3_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_3_tile_v_0_MPORT_3_en = handshaked & _GEN_1317;
  assign rf_matrix_b_3_tile_v_0_MPORT_3_addr = 8'h4e;
  assign rf_matrix_b_3_tile_v_0_MPORT_3_data = rf[rf_matrix_b_3_tile_v_0_MPORT_3_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_3_tile_v_3_MPORT_3_en = handshaked & _GEN_1317;
  assign rf_matrix_c_3_tile_v_3_MPORT_3_addr = 8'ha3;
  assign rf_matrix_c_3_tile_v_3_MPORT_3_data = rf[rf_matrix_c_3_tile_v_3_MPORT_3_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_3_tile_v_2_MPORT_3_en = handshaked & _GEN_1317;
  assign rf_matrix_c_3_tile_v_2_MPORT_3_addr = 8'ha7;
  assign rf_matrix_c_3_tile_v_2_MPORT_3_data = rf[rf_matrix_c_3_tile_v_2_MPORT_3_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_3_tile_v_1_MPORT_3_en = handshaked & _GEN_1317;
  assign rf_matrix_c_3_tile_v_1_MPORT_3_addr = 8'hab;
  assign rf_matrix_c_3_tile_v_1_MPORT_3_data = rf[rf_matrix_c_3_tile_v_1_MPORT_3_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_3_tile_v_0_MPORT_3_en = handshaked & _GEN_1317;
  assign rf_matrix_c_3_tile_v_0_MPORT_3_addr = 8'haf;
  assign rf_matrix_c_3_tile_v_0_MPORT_3_data = rf[rf_matrix_c_3_tile_v_0_MPORT_3_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_1_MPORT_76_en = handshaked & _GEN_1331;
  assign rf_a_tile_v_1_MPORT_76_addr = 8'h20;
  assign rf_a_tile_v_1_MPORT_76_data = rf[rf_a_tile_v_1_MPORT_76_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_0_MPORT_76_en = handshaked & _GEN_1331;
  assign rf_a_tile_v_0_MPORT_76_addr = 8'h24;
  assign rf_a_tile_v_0_MPORT_76_data = rf[rf_a_tile_v_0_MPORT_76_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_3_tile_v_3_MPORT_4_en = handshaked & _GEN_1331;
  assign rf_matrix_b_3_tile_v_3_MPORT_4_addr = 8'h42;
  assign rf_matrix_b_3_tile_v_3_MPORT_4_data = rf[rf_matrix_b_3_tile_v_3_MPORT_4_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_3_tile_v_2_MPORT_4_en = handshaked & _GEN_1331;
  assign rf_matrix_b_3_tile_v_2_MPORT_4_addr = 8'h46;
  assign rf_matrix_b_3_tile_v_2_MPORT_4_data = rf[rf_matrix_b_3_tile_v_2_MPORT_4_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_3_tile_v_1_MPORT_4_en = handshaked & _GEN_1331;
  assign rf_matrix_b_3_tile_v_1_MPORT_4_addr = 8'h4a;
  assign rf_matrix_b_3_tile_v_1_MPORT_4_data = rf[rf_matrix_b_3_tile_v_1_MPORT_4_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_3_tile_v_0_MPORT_4_en = handshaked & _GEN_1331;
  assign rf_matrix_b_3_tile_v_0_MPORT_4_addr = 8'h4e;
  assign rf_matrix_b_3_tile_v_0_MPORT_4_data = rf[rf_matrix_b_3_tile_v_0_MPORT_4_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_3_tile_v_3_MPORT_4_en = handshaked & _GEN_1331;
  assign rf_matrix_c_3_tile_v_3_MPORT_4_addr = 8'hc6;
  assign rf_matrix_c_3_tile_v_3_MPORT_4_data = rf[rf_matrix_c_3_tile_v_3_MPORT_4_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_3_tile_v_2_MPORT_4_en = handshaked & _GEN_1331;
  assign rf_matrix_c_3_tile_v_2_MPORT_4_addr = 8'hc7;
  assign rf_matrix_c_3_tile_v_2_MPORT_4_data = rf[rf_matrix_c_3_tile_v_2_MPORT_4_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_3_tile_v_1_MPORT_4_en = handshaked & _GEN_1331;
  assign rf_matrix_c_3_tile_v_1_MPORT_4_addr = 8'hce;
  assign rf_matrix_c_3_tile_v_1_MPORT_4_data = rf[rf_matrix_c_3_tile_v_1_MPORT_4_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_3_tile_v_0_MPORT_4_en = handshaked & _GEN_1331;
  assign rf_matrix_c_3_tile_v_0_MPORT_4_addr = 8'hcf;
  assign rf_matrix_c_3_tile_v_0_MPORT_4_data = rf[rf_matrix_c_3_tile_v_0_MPORT_4_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_1_MPORT_77_en = handshaked & _GEN_1343;
  assign rf_a_tile_v_1_MPORT_77_addr = 8'h28;
  assign rf_a_tile_v_1_MPORT_77_data = rf[rf_a_tile_v_1_MPORT_77_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_0_MPORT_77_en = handshaked & _GEN_1343;
  assign rf_a_tile_v_0_MPORT_77_addr = 8'h2c;
  assign rf_a_tile_v_0_MPORT_77_data = rf[rf_a_tile_v_0_MPORT_77_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_3_tile_v_3_MPORT_5_en = handshaked & _GEN_1343;
  assign rf_matrix_b_3_tile_v_3_MPORT_5_addr = 8'h42;
  assign rf_matrix_b_3_tile_v_3_MPORT_5_data = rf[rf_matrix_b_3_tile_v_3_MPORT_5_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_3_tile_v_2_MPORT_5_en = handshaked & _GEN_1343;
  assign rf_matrix_b_3_tile_v_2_MPORT_5_addr = 8'h46;
  assign rf_matrix_b_3_tile_v_2_MPORT_5_data = rf[rf_matrix_b_3_tile_v_2_MPORT_5_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_3_tile_v_1_MPORT_5_en = handshaked & _GEN_1343;
  assign rf_matrix_b_3_tile_v_1_MPORT_5_addr = 8'h4a;
  assign rf_matrix_b_3_tile_v_1_MPORT_5_data = rf[rf_matrix_b_3_tile_v_1_MPORT_5_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_3_tile_v_0_MPORT_5_en = handshaked & _GEN_1343;
  assign rf_matrix_b_3_tile_v_0_MPORT_5_addr = 8'h4e;
  assign rf_matrix_b_3_tile_v_0_MPORT_5_data = rf[rf_matrix_b_3_tile_v_0_MPORT_5_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_3_tile_v_3_MPORT_5_en = handshaked & _GEN_1343;
  assign rf_matrix_c_3_tile_v_3_MPORT_5_addr = 8'hd6;
  assign rf_matrix_c_3_tile_v_3_MPORT_5_data = rf[rf_matrix_c_3_tile_v_3_MPORT_5_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_3_tile_v_2_MPORT_5_en = handshaked & _GEN_1343;
  assign rf_matrix_c_3_tile_v_2_MPORT_5_addr = 8'hd7;
  assign rf_matrix_c_3_tile_v_2_MPORT_5_data = rf[rf_matrix_c_3_tile_v_2_MPORT_5_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_3_tile_v_1_MPORT_5_en = handshaked & _GEN_1343;
  assign rf_matrix_c_3_tile_v_1_MPORT_5_addr = 8'hde;
  assign rf_matrix_c_3_tile_v_1_MPORT_5_data = rf[rf_matrix_c_3_tile_v_1_MPORT_5_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_3_tile_v_0_MPORT_5_en = handshaked & _GEN_1343;
  assign rf_matrix_c_3_tile_v_0_MPORT_5_addr = 8'hdf;
  assign rf_matrix_c_3_tile_v_0_MPORT_5_data = rf[rf_matrix_c_3_tile_v_0_MPORT_5_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_1_MPORT_78_en = handshaked & _GEN_1355;
  assign rf_a_tile_v_1_MPORT_78_addr = 8'h21;
  assign rf_a_tile_v_1_MPORT_78_data = rf[rf_a_tile_v_1_MPORT_78_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_0_MPORT_78_en = handshaked & _GEN_1355;
  assign rf_a_tile_v_0_MPORT_78_addr = 8'h25;
  assign rf_a_tile_v_0_MPORT_78_data = rf[rf_a_tile_v_0_MPORT_78_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_3_tile_v_3_MPORT_6_en = handshaked & _GEN_1355;
  assign rf_matrix_b_3_tile_v_3_MPORT_6_addr = 8'h52;
  assign rf_matrix_b_3_tile_v_3_MPORT_6_data = rf[rf_matrix_b_3_tile_v_3_MPORT_6_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_3_tile_v_2_MPORT_6_en = handshaked & _GEN_1355;
  assign rf_matrix_b_3_tile_v_2_MPORT_6_addr = 8'h56;
  assign rf_matrix_b_3_tile_v_2_MPORT_6_data = rf[rf_matrix_b_3_tile_v_2_MPORT_6_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_3_tile_v_1_MPORT_6_en = handshaked & _GEN_1355;
  assign rf_matrix_b_3_tile_v_1_MPORT_6_addr = 8'h5a;
  assign rf_matrix_b_3_tile_v_1_MPORT_6_data = rf[rf_matrix_b_3_tile_v_1_MPORT_6_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_3_tile_v_0_MPORT_6_en = handshaked & _GEN_1355;
  assign rf_matrix_b_3_tile_v_0_MPORT_6_addr = 8'h5e;
  assign rf_matrix_b_3_tile_v_0_MPORT_6_data = rf[rf_matrix_b_3_tile_v_0_MPORT_6_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_3_tile_v_3_MPORT_6_en = handshaked & _GEN_1355;
  assign rf_matrix_c_3_tile_v_3_MPORT_6_addr = 8'hc4;
  assign rf_matrix_c_3_tile_v_3_MPORT_6_data = rf[rf_matrix_c_3_tile_v_3_MPORT_6_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_3_tile_v_2_MPORT_6_en = handshaked & _GEN_1355;
  assign rf_matrix_c_3_tile_v_2_MPORT_6_addr = 8'hc5;
  assign rf_matrix_c_3_tile_v_2_MPORT_6_data = rf[rf_matrix_c_3_tile_v_2_MPORT_6_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_3_tile_v_1_MPORT_6_en = handshaked & _GEN_1355;
  assign rf_matrix_c_3_tile_v_1_MPORT_6_addr = 8'hcc;
  assign rf_matrix_c_3_tile_v_1_MPORT_6_data = rf[rf_matrix_c_3_tile_v_1_MPORT_6_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_3_tile_v_0_MPORT_6_en = handshaked & _GEN_1355;
  assign rf_matrix_c_3_tile_v_0_MPORT_6_addr = 8'hcd;
  assign rf_matrix_c_3_tile_v_0_MPORT_6_data = rf[rf_matrix_c_3_tile_v_0_MPORT_6_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_3_MPORT_26_en = handshaked & _GEN_1367;
  assign rf_a_tile_v_3_MPORT_26_addr = 8'h21;
  assign rf_a_tile_v_3_MPORT_26_data = rf[rf_a_tile_v_3_MPORT_26_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_2_MPORT_26_en = handshaked & _GEN_1367;
  assign rf_a_tile_v_2_MPORT_26_addr = 8'h25;
  assign rf_a_tile_v_2_MPORT_26_data = rf[rf_a_tile_v_2_MPORT_26_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_1_MPORT_79_en = handshaked & _GEN_1367;
  assign rf_a_tile_v_1_MPORT_79_addr = 8'h29;
  assign rf_a_tile_v_1_MPORT_79_data = rf[rf_a_tile_v_1_MPORT_79_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_0_MPORT_79_en = handshaked & _GEN_1367;
  assign rf_a_tile_v_0_MPORT_79_addr = 8'h2d;
  assign rf_a_tile_v_0_MPORT_79_data = rf[rf_a_tile_v_0_MPORT_79_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_3_tile_v_3_MPORT_7_en = handshaked & _GEN_1367;
  assign rf_matrix_b_3_tile_v_3_MPORT_7_addr = 8'h52;
  assign rf_matrix_b_3_tile_v_3_MPORT_7_data = rf[rf_matrix_b_3_tile_v_3_MPORT_7_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_3_tile_v_2_MPORT_7_en = handshaked & _GEN_1367;
  assign rf_matrix_b_3_tile_v_2_MPORT_7_addr = 8'h56;
  assign rf_matrix_b_3_tile_v_2_MPORT_7_data = rf[rf_matrix_b_3_tile_v_2_MPORT_7_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_3_tile_v_1_MPORT_7_en = handshaked & _GEN_1367;
  assign rf_matrix_b_3_tile_v_1_MPORT_7_addr = 8'h5a;
  assign rf_matrix_b_3_tile_v_1_MPORT_7_data = rf[rf_matrix_b_3_tile_v_1_MPORT_7_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_3_tile_v_0_MPORT_7_en = handshaked & _GEN_1367;
  assign rf_matrix_b_3_tile_v_0_MPORT_7_addr = 8'h5e;
  assign rf_matrix_b_3_tile_v_0_MPORT_7_data = rf[rf_matrix_b_3_tile_v_0_MPORT_7_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_3_tile_v_3_MPORT_7_en = handshaked & _GEN_1367;
  assign rf_matrix_c_3_tile_v_3_MPORT_7_addr = 8'ha2;
  assign rf_matrix_c_3_tile_v_3_MPORT_7_data = rf[rf_matrix_c_3_tile_v_3_MPORT_7_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_3_tile_v_2_MPORT_7_en = handshaked & _GEN_1367;
  assign rf_matrix_c_3_tile_v_2_MPORT_7_addr = 8'ha6;
  assign rf_matrix_c_3_tile_v_2_MPORT_7_data = rf[rf_matrix_c_3_tile_v_2_MPORT_7_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_3_tile_v_1_MPORT_7_en = handshaked & _GEN_1367;
  assign rf_matrix_c_3_tile_v_1_MPORT_7_addr = 8'haa;
  assign rf_matrix_c_3_tile_v_1_MPORT_7_data = rf[rf_matrix_c_3_tile_v_1_MPORT_7_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_3_tile_v_0_MPORT_7_en = handshaked & _GEN_1367;
  assign rf_matrix_c_3_tile_v_0_MPORT_7_addr = 8'hae;
  assign rf_matrix_c_3_tile_v_0_MPORT_7_data = rf[rf_matrix_c_3_tile_v_0_MPORT_7_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_1_MPORT_80_en = handshaked & _GEN_1381;
  assign rf_a_tile_v_1_MPORT_80_addr = 8'h29;
  assign rf_a_tile_v_1_MPORT_80_data = rf[rf_a_tile_v_1_MPORT_80_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_0_MPORT_80_en = handshaked & _GEN_1381;
  assign rf_a_tile_v_0_MPORT_80_addr = 8'h2d;
  assign rf_a_tile_v_0_MPORT_80_data = rf[rf_a_tile_v_0_MPORT_80_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_3_tile_v_3_MPORT_8_en = handshaked & _GEN_1381;
  assign rf_matrix_b_3_tile_v_3_MPORT_8_addr = 8'h52;
  assign rf_matrix_b_3_tile_v_3_MPORT_8_data = rf[rf_matrix_b_3_tile_v_3_MPORT_8_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_3_tile_v_2_MPORT_8_en = handshaked & _GEN_1381;
  assign rf_matrix_b_3_tile_v_2_MPORT_8_addr = 8'h56;
  assign rf_matrix_b_3_tile_v_2_MPORT_8_data = rf[rf_matrix_b_3_tile_v_2_MPORT_8_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_3_tile_v_1_MPORT_8_en = handshaked & _GEN_1381;
  assign rf_matrix_b_3_tile_v_1_MPORT_8_addr = 8'h5a;
  assign rf_matrix_b_3_tile_v_1_MPORT_8_data = rf[rf_matrix_b_3_tile_v_1_MPORT_8_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_3_tile_v_0_MPORT_8_en = handshaked & _GEN_1381;
  assign rf_matrix_b_3_tile_v_0_MPORT_8_addr = 8'h5e;
  assign rf_matrix_b_3_tile_v_0_MPORT_8_data = rf[rf_matrix_b_3_tile_v_0_MPORT_8_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_3_tile_v_3_MPORT_8_en = handshaked & _GEN_1381;
  assign rf_matrix_c_3_tile_v_3_MPORT_8_addr = 8'hd4;
  assign rf_matrix_c_3_tile_v_3_MPORT_8_data = rf[rf_matrix_c_3_tile_v_3_MPORT_8_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_3_tile_v_2_MPORT_8_en = handshaked & _GEN_1381;
  assign rf_matrix_c_3_tile_v_2_MPORT_8_addr = 8'hd5;
  assign rf_matrix_c_3_tile_v_2_MPORT_8_data = rf[rf_matrix_c_3_tile_v_2_MPORT_8_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_3_tile_v_1_MPORT_8_en = handshaked & _GEN_1381;
  assign rf_matrix_c_3_tile_v_1_MPORT_8_addr = 8'hdc;
  assign rf_matrix_c_3_tile_v_1_MPORT_8_data = rf[rf_matrix_c_3_tile_v_1_MPORT_8_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_3_tile_v_0_MPORT_8_en = handshaked & _GEN_1381;
  assign rf_matrix_c_3_tile_v_0_MPORT_8_addr = 8'hdd;
  assign rf_matrix_c_3_tile_v_0_MPORT_8_data = rf[rf_matrix_c_3_tile_v_0_MPORT_8_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_3_MPORT_27_en = handshaked & _GEN_1393;
  assign rf_a_tile_v_3_MPORT_27_addr = 8'h21;
  assign rf_a_tile_v_3_MPORT_27_data = rf[rf_a_tile_v_3_MPORT_27_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_2_MPORT_27_en = handshaked & _GEN_1393;
  assign rf_a_tile_v_2_MPORT_27_addr = 8'h25;
  assign rf_a_tile_v_2_MPORT_27_data = rf[rf_a_tile_v_2_MPORT_27_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_1_MPORT_81_en = handshaked & _GEN_1393;
  assign rf_a_tile_v_1_MPORT_81_addr = 8'h29;
  assign rf_a_tile_v_1_MPORT_81_data = rf[rf_a_tile_v_1_MPORT_81_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_0_MPORT_81_en = handshaked & _GEN_1393;
  assign rf_a_tile_v_0_MPORT_81_addr = 8'h2d;
  assign rf_a_tile_v_0_MPORT_81_data = rf[rf_a_tile_v_0_MPORT_81_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_3_tile_v_3_MPORT_9_en = handshaked & _GEN_1393;
  assign rf_matrix_b_3_tile_v_3_MPORT_9_addr = 8'h52;
  assign rf_matrix_b_3_tile_v_3_MPORT_9_data = rf[rf_matrix_b_3_tile_v_3_MPORT_9_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_3_tile_v_2_MPORT_9_en = handshaked & _GEN_1393;
  assign rf_matrix_b_3_tile_v_2_MPORT_9_addr = 8'h56;
  assign rf_matrix_b_3_tile_v_2_MPORT_9_data = rf[rf_matrix_b_3_tile_v_2_MPORT_9_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_3_tile_v_1_MPORT_9_en = handshaked & _GEN_1393;
  assign rf_matrix_b_3_tile_v_1_MPORT_9_addr = 8'h5a;
  assign rf_matrix_b_3_tile_v_1_MPORT_9_data = rf[rf_matrix_b_3_tile_v_1_MPORT_9_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_3_tile_v_0_MPORT_9_en = handshaked & _GEN_1393;
  assign rf_matrix_b_3_tile_v_0_MPORT_9_addr = 8'h5e;
  assign rf_matrix_b_3_tile_v_0_MPORT_9_data = rf[rf_matrix_b_3_tile_v_0_MPORT_9_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_3_tile_v_3_MPORT_9_en = handshaked & _GEN_1393;
  assign rf_matrix_c_3_tile_v_3_MPORT_9_addr = 8'ha3;
  assign rf_matrix_c_3_tile_v_3_MPORT_9_data = rf[rf_matrix_c_3_tile_v_3_MPORT_9_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_3_tile_v_2_MPORT_9_en = handshaked & _GEN_1393;
  assign rf_matrix_c_3_tile_v_2_MPORT_9_addr = 8'ha7;
  assign rf_matrix_c_3_tile_v_2_MPORT_9_data = rf[rf_matrix_c_3_tile_v_2_MPORT_9_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_3_tile_v_1_MPORT_9_en = handshaked & _GEN_1393;
  assign rf_matrix_c_3_tile_v_1_MPORT_9_addr = 8'hab;
  assign rf_matrix_c_3_tile_v_1_MPORT_9_data = rf[rf_matrix_c_3_tile_v_1_MPORT_9_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_3_tile_v_0_MPORT_9_en = handshaked & _GEN_1393;
  assign rf_matrix_c_3_tile_v_0_MPORT_9_addr = 8'haf;
  assign rf_matrix_c_3_tile_v_0_MPORT_9_data = rf[rf_matrix_c_3_tile_v_0_MPORT_9_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_1_MPORT_82_en = handshaked & _GEN_1407;
  assign rf_a_tile_v_1_MPORT_82_addr = 8'h21;
  assign rf_a_tile_v_1_MPORT_82_data = rf[rf_a_tile_v_1_MPORT_82_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_0_MPORT_82_en = handshaked & _GEN_1407;
  assign rf_a_tile_v_0_MPORT_82_addr = 8'h25;
  assign rf_a_tile_v_0_MPORT_82_data = rf[rf_a_tile_v_0_MPORT_82_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_3_tile_v_3_MPORT_10_en = handshaked & _GEN_1407;
  assign rf_matrix_b_3_tile_v_3_MPORT_10_addr = 8'h52;
  assign rf_matrix_b_3_tile_v_3_MPORT_10_data = rf[rf_matrix_b_3_tile_v_3_MPORT_10_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_3_tile_v_2_MPORT_10_en = handshaked & _GEN_1407;
  assign rf_matrix_b_3_tile_v_2_MPORT_10_addr = 8'h56;
  assign rf_matrix_b_3_tile_v_2_MPORT_10_data = rf[rf_matrix_b_3_tile_v_2_MPORT_10_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_3_tile_v_1_MPORT_10_en = handshaked & _GEN_1407;
  assign rf_matrix_b_3_tile_v_1_MPORT_10_addr = 8'h5a;
  assign rf_matrix_b_3_tile_v_1_MPORT_10_data = rf[rf_matrix_b_3_tile_v_1_MPORT_10_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_3_tile_v_0_MPORT_10_en = handshaked & _GEN_1407;
  assign rf_matrix_b_3_tile_v_0_MPORT_10_addr = 8'h5e;
  assign rf_matrix_b_3_tile_v_0_MPORT_10_data = rf[rf_matrix_b_3_tile_v_0_MPORT_10_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_3_tile_v_3_MPORT_10_en = handshaked & _GEN_1407;
  assign rf_matrix_c_3_tile_v_3_MPORT_10_addr = 8'hc6;
  assign rf_matrix_c_3_tile_v_3_MPORT_10_data = rf[rf_matrix_c_3_tile_v_3_MPORT_10_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_3_tile_v_2_MPORT_10_en = handshaked & _GEN_1407;
  assign rf_matrix_c_3_tile_v_2_MPORT_10_addr = 8'hc7;
  assign rf_matrix_c_3_tile_v_2_MPORT_10_data = rf[rf_matrix_c_3_tile_v_2_MPORT_10_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_3_tile_v_1_MPORT_10_en = handshaked & _GEN_1407;
  assign rf_matrix_c_3_tile_v_1_MPORT_10_addr = 8'hce;
  assign rf_matrix_c_3_tile_v_1_MPORT_10_data = rf[rf_matrix_c_3_tile_v_1_MPORT_10_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_3_tile_v_0_MPORT_10_en = handshaked & _GEN_1407;
  assign rf_matrix_c_3_tile_v_0_MPORT_10_addr = 8'hcf;
  assign rf_matrix_c_3_tile_v_0_MPORT_10_data = rf[rf_matrix_c_3_tile_v_0_MPORT_10_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_1_MPORT_83_en = handshaked & _GEN_1419;
  assign rf_a_tile_v_1_MPORT_83_addr = 8'h29;
  assign rf_a_tile_v_1_MPORT_83_data = rf[rf_a_tile_v_1_MPORT_83_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_0_MPORT_83_en = handshaked & _GEN_1419;
  assign rf_a_tile_v_0_MPORT_83_addr = 8'h2d;
  assign rf_a_tile_v_0_MPORT_83_data = rf[rf_a_tile_v_0_MPORT_83_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_3_tile_v_3_MPORT_11_en = handshaked & _GEN_1419;
  assign rf_matrix_b_3_tile_v_3_MPORT_11_addr = 8'h52;
  assign rf_matrix_b_3_tile_v_3_MPORT_11_data = rf[rf_matrix_b_3_tile_v_3_MPORT_11_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_3_tile_v_2_MPORT_11_en = handshaked & _GEN_1419;
  assign rf_matrix_b_3_tile_v_2_MPORT_11_addr = 8'h56;
  assign rf_matrix_b_3_tile_v_2_MPORT_11_data = rf[rf_matrix_b_3_tile_v_2_MPORT_11_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_3_tile_v_1_MPORT_11_en = handshaked & _GEN_1419;
  assign rf_matrix_b_3_tile_v_1_MPORT_11_addr = 8'h5a;
  assign rf_matrix_b_3_tile_v_1_MPORT_11_data = rf[rf_matrix_b_3_tile_v_1_MPORT_11_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_3_tile_v_0_MPORT_11_en = handshaked & _GEN_1419;
  assign rf_matrix_b_3_tile_v_0_MPORT_11_addr = 8'h5e;
  assign rf_matrix_b_3_tile_v_0_MPORT_11_data = rf[rf_matrix_b_3_tile_v_0_MPORT_11_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_3_tile_v_3_MPORT_11_en = handshaked & _GEN_1419;
  assign rf_matrix_c_3_tile_v_3_MPORT_11_addr = 8'hd6;
  assign rf_matrix_c_3_tile_v_3_MPORT_11_data = rf[rf_matrix_c_3_tile_v_3_MPORT_11_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_3_tile_v_2_MPORT_11_en = handshaked & _GEN_1419;
  assign rf_matrix_c_3_tile_v_2_MPORT_11_addr = 8'hd7;
  assign rf_matrix_c_3_tile_v_2_MPORT_11_data = rf[rf_matrix_c_3_tile_v_2_MPORT_11_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_3_tile_v_1_MPORT_11_en = handshaked & _GEN_1419;
  assign rf_matrix_c_3_tile_v_1_MPORT_11_addr = 8'hde;
  assign rf_matrix_c_3_tile_v_1_MPORT_11_data = rf[rf_matrix_c_3_tile_v_1_MPORT_11_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_3_tile_v_0_MPORT_11_en = handshaked & _GEN_1419;
  assign rf_matrix_c_3_tile_v_0_MPORT_11_addr = 8'hdf;
  assign rf_matrix_c_3_tile_v_0_MPORT_11_data = rf[rf_matrix_c_3_tile_v_0_MPORT_11_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_1_MPORT_84_en = handshaked & _GEN_1431;
  assign rf_a_tile_v_1_MPORT_84_addr = 8'h22;
  assign rf_a_tile_v_1_MPORT_84_data = rf[rf_a_tile_v_1_MPORT_84_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_0_MPORT_84_en = handshaked & _GEN_1431;
  assign rf_a_tile_v_0_MPORT_84_addr = 8'h26;
  assign rf_a_tile_v_0_MPORT_84_data = rf[rf_a_tile_v_0_MPORT_84_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_3_tile_v_3_MPORT_12_en = handshaked & _GEN_1431;
  assign rf_matrix_b_3_tile_v_3_MPORT_12_addr = 8'h62;
  assign rf_matrix_b_3_tile_v_3_MPORT_12_data = rf[rf_matrix_b_3_tile_v_3_MPORT_12_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_3_tile_v_2_MPORT_12_en = handshaked & _GEN_1431;
  assign rf_matrix_b_3_tile_v_2_MPORT_12_addr = 8'h66;
  assign rf_matrix_b_3_tile_v_2_MPORT_12_data = rf[rf_matrix_b_3_tile_v_2_MPORT_12_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_3_tile_v_1_MPORT_12_en = handshaked & _GEN_1431;
  assign rf_matrix_b_3_tile_v_1_MPORT_12_addr = 8'h6a;
  assign rf_matrix_b_3_tile_v_1_MPORT_12_data = rf[rf_matrix_b_3_tile_v_1_MPORT_12_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_3_tile_v_0_MPORT_12_en = handshaked & _GEN_1431;
  assign rf_matrix_b_3_tile_v_0_MPORT_12_addr = 8'h6e;
  assign rf_matrix_b_3_tile_v_0_MPORT_12_data = rf[rf_matrix_b_3_tile_v_0_MPORT_12_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_3_tile_v_3_MPORT_12_en = handshaked & _GEN_1431;
  assign rf_matrix_c_3_tile_v_3_MPORT_12_addr = 8'hc4;
  assign rf_matrix_c_3_tile_v_3_MPORT_12_data = rf[rf_matrix_c_3_tile_v_3_MPORT_12_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_3_tile_v_2_MPORT_12_en = handshaked & _GEN_1431;
  assign rf_matrix_c_3_tile_v_2_MPORT_12_addr = 8'hc5;
  assign rf_matrix_c_3_tile_v_2_MPORT_12_data = rf[rf_matrix_c_3_tile_v_2_MPORT_12_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_3_tile_v_1_MPORT_12_en = handshaked & _GEN_1431;
  assign rf_matrix_c_3_tile_v_1_MPORT_12_addr = 8'hcc;
  assign rf_matrix_c_3_tile_v_1_MPORT_12_data = rf[rf_matrix_c_3_tile_v_1_MPORT_12_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_3_tile_v_0_MPORT_12_en = handshaked & _GEN_1431;
  assign rf_matrix_c_3_tile_v_0_MPORT_12_addr = 8'hcd;
  assign rf_matrix_c_3_tile_v_0_MPORT_12_data = rf[rf_matrix_c_3_tile_v_0_MPORT_12_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_3_MPORT_28_en = handshaked & _GEN_1443;
  assign rf_a_tile_v_3_MPORT_28_addr = 8'h22;
  assign rf_a_tile_v_3_MPORT_28_data = rf[rf_a_tile_v_3_MPORT_28_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_2_MPORT_28_en = handshaked & _GEN_1443;
  assign rf_a_tile_v_2_MPORT_28_addr = 8'h26;
  assign rf_a_tile_v_2_MPORT_28_data = rf[rf_a_tile_v_2_MPORT_28_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_1_MPORT_85_en = handshaked & _GEN_1443;
  assign rf_a_tile_v_1_MPORT_85_addr = 8'h2a;
  assign rf_a_tile_v_1_MPORT_85_data = rf[rf_a_tile_v_1_MPORT_85_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_0_MPORT_85_en = handshaked & _GEN_1443;
  assign rf_a_tile_v_0_MPORT_85_addr = 8'h2e;
  assign rf_a_tile_v_0_MPORT_85_data = rf[rf_a_tile_v_0_MPORT_85_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_3_tile_v_3_MPORT_13_en = handshaked & _GEN_1443;
  assign rf_matrix_b_3_tile_v_3_MPORT_13_addr = 8'h62;
  assign rf_matrix_b_3_tile_v_3_MPORT_13_data = rf[rf_matrix_b_3_tile_v_3_MPORT_13_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_3_tile_v_2_MPORT_13_en = handshaked & _GEN_1443;
  assign rf_matrix_b_3_tile_v_2_MPORT_13_addr = 8'h66;
  assign rf_matrix_b_3_tile_v_2_MPORT_13_data = rf[rf_matrix_b_3_tile_v_2_MPORT_13_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_3_tile_v_1_MPORT_13_en = handshaked & _GEN_1443;
  assign rf_matrix_b_3_tile_v_1_MPORT_13_addr = 8'h6a;
  assign rf_matrix_b_3_tile_v_1_MPORT_13_data = rf[rf_matrix_b_3_tile_v_1_MPORT_13_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_3_tile_v_0_MPORT_13_en = handshaked & _GEN_1443;
  assign rf_matrix_b_3_tile_v_0_MPORT_13_addr = 8'h6e;
  assign rf_matrix_b_3_tile_v_0_MPORT_13_data = rf[rf_matrix_b_3_tile_v_0_MPORT_13_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_3_tile_v_3_MPORT_13_en = handshaked & _GEN_1443;
  assign rf_matrix_c_3_tile_v_3_MPORT_13_addr = 8'ha2;
  assign rf_matrix_c_3_tile_v_3_MPORT_13_data = rf[rf_matrix_c_3_tile_v_3_MPORT_13_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_3_tile_v_2_MPORT_13_en = handshaked & _GEN_1443;
  assign rf_matrix_c_3_tile_v_2_MPORT_13_addr = 8'ha6;
  assign rf_matrix_c_3_tile_v_2_MPORT_13_data = rf[rf_matrix_c_3_tile_v_2_MPORT_13_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_3_tile_v_1_MPORT_13_en = handshaked & _GEN_1443;
  assign rf_matrix_c_3_tile_v_1_MPORT_13_addr = 8'haa;
  assign rf_matrix_c_3_tile_v_1_MPORT_13_data = rf[rf_matrix_c_3_tile_v_1_MPORT_13_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_3_tile_v_0_MPORT_13_en = handshaked & _GEN_1443;
  assign rf_matrix_c_3_tile_v_0_MPORT_13_addr = 8'hae;
  assign rf_matrix_c_3_tile_v_0_MPORT_13_data = rf[rf_matrix_c_3_tile_v_0_MPORT_13_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_1_MPORT_86_en = handshaked & _GEN_1457;
  assign rf_a_tile_v_1_MPORT_86_addr = 8'h2a;
  assign rf_a_tile_v_1_MPORT_86_data = rf[rf_a_tile_v_1_MPORT_86_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_0_MPORT_86_en = handshaked & _GEN_1457;
  assign rf_a_tile_v_0_MPORT_86_addr = 8'h2e;
  assign rf_a_tile_v_0_MPORT_86_data = rf[rf_a_tile_v_0_MPORT_86_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_3_tile_v_3_MPORT_14_en = handshaked & _GEN_1457;
  assign rf_matrix_b_3_tile_v_3_MPORT_14_addr = 8'h62;
  assign rf_matrix_b_3_tile_v_3_MPORT_14_data = rf[rf_matrix_b_3_tile_v_3_MPORT_14_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_3_tile_v_2_MPORT_14_en = handshaked & _GEN_1457;
  assign rf_matrix_b_3_tile_v_2_MPORT_14_addr = 8'h66;
  assign rf_matrix_b_3_tile_v_2_MPORT_14_data = rf[rf_matrix_b_3_tile_v_2_MPORT_14_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_3_tile_v_1_MPORT_14_en = handshaked & _GEN_1457;
  assign rf_matrix_b_3_tile_v_1_MPORT_14_addr = 8'h6a;
  assign rf_matrix_b_3_tile_v_1_MPORT_14_data = rf[rf_matrix_b_3_tile_v_1_MPORT_14_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_3_tile_v_0_MPORT_14_en = handshaked & _GEN_1457;
  assign rf_matrix_b_3_tile_v_0_MPORT_14_addr = 8'h6e;
  assign rf_matrix_b_3_tile_v_0_MPORT_14_data = rf[rf_matrix_b_3_tile_v_0_MPORT_14_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_3_tile_v_3_MPORT_14_en = handshaked & _GEN_1457;
  assign rf_matrix_c_3_tile_v_3_MPORT_14_addr = 8'hd4;
  assign rf_matrix_c_3_tile_v_3_MPORT_14_data = rf[rf_matrix_c_3_tile_v_3_MPORT_14_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_3_tile_v_2_MPORT_14_en = handshaked & _GEN_1457;
  assign rf_matrix_c_3_tile_v_2_MPORT_14_addr = 8'hd5;
  assign rf_matrix_c_3_tile_v_2_MPORT_14_data = rf[rf_matrix_c_3_tile_v_2_MPORT_14_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_3_tile_v_1_MPORT_14_en = handshaked & _GEN_1457;
  assign rf_matrix_c_3_tile_v_1_MPORT_14_addr = 8'hdc;
  assign rf_matrix_c_3_tile_v_1_MPORT_14_data = rf[rf_matrix_c_3_tile_v_1_MPORT_14_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_3_tile_v_0_MPORT_14_en = handshaked & _GEN_1457;
  assign rf_matrix_c_3_tile_v_0_MPORT_14_addr = 8'hdd;
  assign rf_matrix_c_3_tile_v_0_MPORT_14_data = rf[rf_matrix_c_3_tile_v_0_MPORT_14_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_3_MPORT_29_en = handshaked & _GEN_1469;
  assign rf_a_tile_v_3_MPORT_29_addr = 8'h22;
  assign rf_a_tile_v_3_MPORT_29_data = rf[rf_a_tile_v_3_MPORT_29_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_2_MPORT_29_en = handshaked & _GEN_1469;
  assign rf_a_tile_v_2_MPORT_29_addr = 8'h26;
  assign rf_a_tile_v_2_MPORT_29_data = rf[rf_a_tile_v_2_MPORT_29_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_1_MPORT_87_en = handshaked & _GEN_1469;
  assign rf_a_tile_v_1_MPORT_87_addr = 8'h2a;
  assign rf_a_tile_v_1_MPORT_87_data = rf[rf_a_tile_v_1_MPORT_87_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_0_MPORT_87_en = handshaked & _GEN_1469;
  assign rf_a_tile_v_0_MPORT_87_addr = 8'h2e;
  assign rf_a_tile_v_0_MPORT_87_data = rf[rf_a_tile_v_0_MPORT_87_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_3_tile_v_3_MPORT_15_en = handshaked & _GEN_1469;
  assign rf_matrix_b_3_tile_v_3_MPORT_15_addr = 8'h62;
  assign rf_matrix_b_3_tile_v_3_MPORT_15_data = rf[rf_matrix_b_3_tile_v_3_MPORT_15_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_3_tile_v_2_MPORT_15_en = handshaked & _GEN_1469;
  assign rf_matrix_b_3_tile_v_2_MPORT_15_addr = 8'h66;
  assign rf_matrix_b_3_tile_v_2_MPORT_15_data = rf[rf_matrix_b_3_tile_v_2_MPORT_15_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_3_tile_v_1_MPORT_15_en = handshaked & _GEN_1469;
  assign rf_matrix_b_3_tile_v_1_MPORT_15_addr = 8'h6a;
  assign rf_matrix_b_3_tile_v_1_MPORT_15_data = rf[rf_matrix_b_3_tile_v_1_MPORT_15_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_3_tile_v_0_MPORT_15_en = handshaked & _GEN_1469;
  assign rf_matrix_b_3_tile_v_0_MPORT_15_addr = 8'h6e;
  assign rf_matrix_b_3_tile_v_0_MPORT_15_data = rf[rf_matrix_b_3_tile_v_0_MPORT_15_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_3_tile_v_3_MPORT_15_en = handshaked & _GEN_1469;
  assign rf_matrix_c_3_tile_v_3_MPORT_15_addr = 8'ha3;
  assign rf_matrix_c_3_tile_v_3_MPORT_15_data = rf[rf_matrix_c_3_tile_v_3_MPORT_15_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_3_tile_v_2_MPORT_15_en = handshaked & _GEN_1469;
  assign rf_matrix_c_3_tile_v_2_MPORT_15_addr = 8'ha7;
  assign rf_matrix_c_3_tile_v_2_MPORT_15_data = rf[rf_matrix_c_3_tile_v_2_MPORT_15_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_3_tile_v_1_MPORT_15_en = handshaked & _GEN_1469;
  assign rf_matrix_c_3_tile_v_1_MPORT_15_addr = 8'hab;
  assign rf_matrix_c_3_tile_v_1_MPORT_15_data = rf[rf_matrix_c_3_tile_v_1_MPORT_15_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_3_tile_v_0_MPORT_15_en = handshaked & _GEN_1469;
  assign rf_matrix_c_3_tile_v_0_MPORT_15_addr = 8'haf;
  assign rf_matrix_c_3_tile_v_0_MPORT_15_data = rf[rf_matrix_c_3_tile_v_0_MPORT_15_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_1_MPORT_88_en = handshaked & _GEN_1483;
  assign rf_a_tile_v_1_MPORT_88_addr = 8'h22;
  assign rf_a_tile_v_1_MPORT_88_data = rf[rf_a_tile_v_1_MPORT_88_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_0_MPORT_88_en = handshaked & _GEN_1483;
  assign rf_a_tile_v_0_MPORT_88_addr = 8'h26;
  assign rf_a_tile_v_0_MPORT_88_data = rf[rf_a_tile_v_0_MPORT_88_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_3_tile_v_3_MPORT_16_en = handshaked & _GEN_1483;
  assign rf_matrix_b_3_tile_v_3_MPORT_16_addr = 8'h62;
  assign rf_matrix_b_3_tile_v_3_MPORT_16_data = rf[rf_matrix_b_3_tile_v_3_MPORT_16_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_3_tile_v_2_MPORT_16_en = handshaked & _GEN_1483;
  assign rf_matrix_b_3_tile_v_2_MPORT_16_addr = 8'h66;
  assign rf_matrix_b_3_tile_v_2_MPORT_16_data = rf[rf_matrix_b_3_tile_v_2_MPORT_16_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_3_tile_v_1_MPORT_16_en = handshaked & _GEN_1483;
  assign rf_matrix_b_3_tile_v_1_MPORT_16_addr = 8'h6a;
  assign rf_matrix_b_3_tile_v_1_MPORT_16_data = rf[rf_matrix_b_3_tile_v_1_MPORT_16_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_3_tile_v_0_MPORT_16_en = handshaked & _GEN_1483;
  assign rf_matrix_b_3_tile_v_0_MPORT_16_addr = 8'h6e;
  assign rf_matrix_b_3_tile_v_0_MPORT_16_data = rf[rf_matrix_b_3_tile_v_0_MPORT_16_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_3_tile_v_3_MPORT_16_en = handshaked & _GEN_1483;
  assign rf_matrix_c_3_tile_v_3_MPORT_16_addr = 8'hc6;
  assign rf_matrix_c_3_tile_v_3_MPORT_16_data = rf[rf_matrix_c_3_tile_v_3_MPORT_16_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_3_tile_v_2_MPORT_16_en = handshaked & _GEN_1483;
  assign rf_matrix_c_3_tile_v_2_MPORT_16_addr = 8'hc7;
  assign rf_matrix_c_3_tile_v_2_MPORT_16_data = rf[rf_matrix_c_3_tile_v_2_MPORT_16_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_3_tile_v_1_MPORT_16_en = handshaked & _GEN_1483;
  assign rf_matrix_c_3_tile_v_1_MPORT_16_addr = 8'hce;
  assign rf_matrix_c_3_tile_v_1_MPORT_16_data = rf[rf_matrix_c_3_tile_v_1_MPORT_16_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_3_tile_v_0_MPORT_16_en = handshaked & _GEN_1483;
  assign rf_matrix_c_3_tile_v_0_MPORT_16_addr = 8'hcf;
  assign rf_matrix_c_3_tile_v_0_MPORT_16_data = rf[rf_matrix_c_3_tile_v_0_MPORT_16_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_1_MPORT_89_en = handshaked & _GEN_1495;
  assign rf_a_tile_v_1_MPORT_89_addr = 8'h2a;
  assign rf_a_tile_v_1_MPORT_89_data = rf[rf_a_tile_v_1_MPORT_89_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_0_MPORT_89_en = handshaked & _GEN_1495;
  assign rf_a_tile_v_0_MPORT_89_addr = 8'h2e;
  assign rf_a_tile_v_0_MPORT_89_data = rf[rf_a_tile_v_0_MPORT_89_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_3_tile_v_3_MPORT_17_en = handshaked & _GEN_1495;
  assign rf_matrix_b_3_tile_v_3_MPORT_17_addr = 8'h62;
  assign rf_matrix_b_3_tile_v_3_MPORT_17_data = rf[rf_matrix_b_3_tile_v_3_MPORT_17_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_3_tile_v_2_MPORT_17_en = handshaked & _GEN_1495;
  assign rf_matrix_b_3_tile_v_2_MPORT_17_addr = 8'h66;
  assign rf_matrix_b_3_tile_v_2_MPORT_17_data = rf[rf_matrix_b_3_tile_v_2_MPORT_17_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_3_tile_v_1_MPORT_17_en = handshaked & _GEN_1495;
  assign rf_matrix_b_3_tile_v_1_MPORT_17_addr = 8'h6a;
  assign rf_matrix_b_3_tile_v_1_MPORT_17_data = rf[rf_matrix_b_3_tile_v_1_MPORT_17_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_3_tile_v_0_MPORT_17_en = handshaked & _GEN_1495;
  assign rf_matrix_b_3_tile_v_0_MPORT_17_addr = 8'h6e;
  assign rf_matrix_b_3_tile_v_0_MPORT_17_data = rf[rf_matrix_b_3_tile_v_0_MPORT_17_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_3_tile_v_3_MPORT_17_en = handshaked & _GEN_1495;
  assign rf_matrix_c_3_tile_v_3_MPORT_17_addr = 8'hd6;
  assign rf_matrix_c_3_tile_v_3_MPORT_17_data = rf[rf_matrix_c_3_tile_v_3_MPORT_17_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_3_tile_v_2_MPORT_17_en = handshaked & _GEN_1495;
  assign rf_matrix_c_3_tile_v_2_MPORT_17_addr = 8'hd7;
  assign rf_matrix_c_3_tile_v_2_MPORT_17_data = rf[rf_matrix_c_3_tile_v_2_MPORT_17_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_3_tile_v_1_MPORT_17_en = handshaked & _GEN_1495;
  assign rf_matrix_c_3_tile_v_1_MPORT_17_addr = 8'hde;
  assign rf_matrix_c_3_tile_v_1_MPORT_17_data = rf[rf_matrix_c_3_tile_v_1_MPORT_17_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_3_tile_v_0_MPORT_17_en = handshaked & _GEN_1495;
  assign rf_matrix_c_3_tile_v_0_MPORT_17_addr = 8'hdf;
  assign rf_matrix_c_3_tile_v_0_MPORT_17_data = rf[rf_matrix_c_3_tile_v_0_MPORT_17_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_1_MPORT_90_en = handshaked & _GEN_1507;
  assign rf_a_tile_v_1_MPORT_90_addr = 8'h23;
  assign rf_a_tile_v_1_MPORT_90_data = rf[rf_a_tile_v_1_MPORT_90_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_0_MPORT_90_en = handshaked & _GEN_1507;
  assign rf_a_tile_v_0_MPORT_90_addr = 8'h27;
  assign rf_a_tile_v_0_MPORT_90_data = rf[rf_a_tile_v_0_MPORT_90_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_3_tile_v_3_MPORT_18_en = handshaked & _GEN_1507;
  assign rf_matrix_b_3_tile_v_3_MPORT_18_addr = 8'h72;
  assign rf_matrix_b_3_tile_v_3_MPORT_18_data = rf[rf_matrix_b_3_tile_v_3_MPORT_18_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_3_tile_v_2_MPORT_18_en = handshaked & _GEN_1507;
  assign rf_matrix_b_3_tile_v_2_MPORT_18_addr = 8'h76;
  assign rf_matrix_b_3_tile_v_2_MPORT_18_data = rf[rf_matrix_b_3_tile_v_2_MPORT_18_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_3_tile_v_1_MPORT_18_en = handshaked & _GEN_1507;
  assign rf_matrix_b_3_tile_v_1_MPORT_18_addr = 8'h7a;
  assign rf_matrix_b_3_tile_v_1_MPORT_18_data = rf[rf_matrix_b_3_tile_v_1_MPORT_18_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_3_tile_v_0_MPORT_18_en = handshaked & _GEN_1507;
  assign rf_matrix_b_3_tile_v_0_MPORT_18_addr = 8'h7e;
  assign rf_matrix_b_3_tile_v_0_MPORT_18_data = rf[rf_matrix_b_3_tile_v_0_MPORT_18_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_3_tile_v_3_MPORT_18_en = handshaked & _GEN_1507;
  assign rf_matrix_c_3_tile_v_3_MPORT_18_addr = 8'hc4;
  assign rf_matrix_c_3_tile_v_3_MPORT_18_data = rf[rf_matrix_c_3_tile_v_3_MPORT_18_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_3_tile_v_2_MPORT_18_en = handshaked & _GEN_1507;
  assign rf_matrix_c_3_tile_v_2_MPORT_18_addr = 8'hc5;
  assign rf_matrix_c_3_tile_v_2_MPORT_18_data = rf[rf_matrix_c_3_tile_v_2_MPORT_18_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_3_tile_v_1_MPORT_18_en = handshaked & _GEN_1507;
  assign rf_matrix_c_3_tile_v_1_MPORT_18_addr = 8'hcc;
  assign rf_matrix_c_3_tile_v_1_MPORT_18_data = rf[rf_matrix_c_3_tile_v_1_MPORT_18_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_3_tile_v_0_MPORT_18_en = handshaked & _GEN_1507;
  assign rf_matrix_c_3_tile_v_0_MPORT_18_addr = 8'hcd;
  assign rf_matrix_c_3_tile_v_0_MPORT_18_data = rf[rf_matrix_c_3_tile_v_0_MPORT_18_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_3_MPORT_30_en = handshaked & _GEN_1519;
  assign rf_a_tile_v_3_MPORT_30_addr = 8'h23;
  assign rf_a_tile_v_3_MPORT_30_data = rf[rf_a_tile_v_3_MPORT_30_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_2_MPORT_30_en = handshaked & _GEN_1519;
  assign rf_a_tile_v_2_MPORT_30_addr = 8'h27;
  assign rf_a_tile_v_2_MPORT_30_data = rf[rf_a_tile_v_2_MPORT_30_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_1_MPORT_91_en = handshaked & _GEN_1519;
  assign rf_a_tile_v_1_MPORT_91_addr = 8'h2b;
  assign rf_a_tile_v_1_MPORT_91_data = rf[rf_a_tile_v_1_MPORT_91_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_0_MPORT_91_en = handshaked & _GEN_1519;
  assign rf_a_tile_v_0_MPORT_91_addr = 8'h2f;
  assign rf_a_tile_v_0_MPORT_91_data = rf[rf_a_tile_v_0_MPORT_91_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_3_tile_v_3_MPORT_19_en = handshaked & _GEN_1519;
  assign rf_matrix_b_3_tile_v_3_MPORT_19_addr = 8'h72;
  assign rf_matrix_b_3_tile_v_3_MPORT_19_data = rf[rf_matrix_b_3_tile_v_3_MPORT_19_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_3_tile_v_2_MPORT_19_en = handshaked & _GEN_1519;
  assign rf_matrix_b_3_tile_v_2_MPORT_19_addr = 8'h76;
  assign rf_matrix_b_3_tile_v_2_MPORT_19_data = rf[rf_matrix_b_3_tile_v_2_MPORT_19_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_3_tile_v_1_MPORT_19_en = handshaked & _GEN_1519;
  assign rf_matrix_b_3_tile_v_1_MPORT_19_addr = 8'h7a;
  assign rf_matrix_b_3_tile_v_1_MPORT_19_data = rf[rf_matrix_b_3_tile_v_1_MPORT_19_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_3_tile_v_0_MPORT_19_en = handshaked & _GEN_1519;
  assign rf_matrix_b_3_tile_v_0_MPORT_19_addr = 8'h7e;
  assign rf_matrix_b_3_tile_v_0_MPORT_19_data = rf[rf_matrix_b_3_tile_v_0_MPORT_19_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_3_tile_v_3_MPORT_19_en = handshaked & _GEN_1519;
  assign rf_matrix_c_3_tile_v_3_MPORT_19_addr = 8'ha2;
  assign rf_matrix_c_3_tile_v_3_MPORT_19_data = rf[rf_matrix_c_3_tile_v_3_MPORT_19_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_3_tile_v_2_MPORT_19_en = handshaked & _GEN_1519;
  assign rf_matrix_c_3_tile_v_2_MPORT_19_addr = 8'ha6;
  assign rf_matrix_c_3_tile_v_2_MPORT_19_data = rf[rf_matrix_c_3_tile_v_2_MPORT_19_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_3_tile_v_1_MPORT_19_en = handshaked & _GEN_1519;
  assign rf_matrix_c_3_tile_v_1_MPORT_19_addr = 8'haa;
  assign rf_matrix_c_3_tile_v_1_MPORT_19_data = rf[rf_matrix_c_3_tile_v_1_MPORT_19_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_3_tile_v_0_MPORT_19_en = handshaked & _GEN_1519;
  assign rf_matrix_c_3_tile_v_0_MPORT_19_addr = 8'hae;
  assign rf_matrix_c_3_tile_v_0_MPORT_19_data = rf[rf_matrix_c_3_tile_v_0_MPORT_19_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_1_MPORT_92_en = handshaked & _GEN_1533;
  assign rf_a_tile_v_1_MPORT_92_addr = 8'h2b;
  assign rf_a_tile_v_1_MPORT_92_data = rf[rf_a_tile_v_1_MPORT_92_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_0_MPORT_92_en = handshaked & _GEN_1533;
  assign rf_a_tile_v_0_MPORT_92_addr = 8'h2f;
  assign rf_a_tile_v_0_MPORT_92_data = rf[rf_a_tile_v_0_MPORT_92_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_3_tile_v_3_MPORT_20_en = handshaked & _GEN_1533;
  assign rf_matrix_b_3_tile_v_3_MPORT_20_addr = 8'h72;
  assign rf_matrix_b_3_tile_v_3_MPORT_20_data = rf[rf_matrix_b_3_tile_v_3_MPORT_20_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_3_tile_v_2_MPORT_20_en = handshaked & _GEN_1533;
  assign rf_matrix_b_3_tile_v_2_MPORT_20_addr = 8'h76;
  assign rf_matrix_b_3_tile_v_2_MPORT_20_data = rf[rf_matrix_b_3_tile_v_2_MPORT_20_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_3_tile_v_1_MPORT_20_en = handshaked & _GEN_1533;
  assign rf_matrix_b_3_tile_v_1_MPORT_20_addr = 8'h7a;
  assign rf_matrix_b_3_tile_v_1_MPORT_20_data = rf[rf_matrix_b_3_tile_v_1_MPORT_20_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_3_tile_v_0_MPORT_20_en = handshaked & _GEN_1533;
  assign rf_matrix_b_3_tile_v_0_MPORT_20_addr = 8'h7e;
  assign rf_matrix_b_3_tile_v_0_MPORT_20_data = rf[rf_matrix_b_3_tile_v_0_MPORT_20_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_3_tile_v_3_MPORT_20_en = handshaked & _GEN_1533;
  assign rf_matrix_c_3_tile_v_3_MPORT_20_addr = 8'hd4;
  assign rf_matrix_c_3_tile_v_3_MPORT_20_data = rf[rf_matrix_c_3_tile_v_3_MPORT_20_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_3_tile_v_2_MPORT_20_en = handshaked & _GEN_1533;
  assign rf_matrix_c_3_tile_v_2_MPORT_20_addr = 8'hd5;
  assign rf_matrix_c_3_tile_v_2_MPORT_20_data = rf[rf_matrix_c_3_tile_v_2_MPORT_20_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_3_tile_v_1_MPORT_20_en = handshaked & _GEN_1533;
  assign rf_matrix_c_3_tile_v_1_MPORT_20_addr = 8'hdc;
  assign rf_matrix_c_3_tile_v_1_MPORT_20_data = rf[rf_matrix_c_3_tile_v_1_MPORT_20_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_3_tile_v_0_MPORT_20_en = handshaked & _GEN_1533;
  assign rf_matrix_c_3_tile_v_0_MPORT_20_addr = 8'hdd;
  assign rf_matrix_c_3_tile_v_0_MPORT_20_data = rf[rf_matrix_c_3_tile_v_0_MPORT_20_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_3_MPORT_31_en = handshaked & _GEN_1545;
  assign rf_a_tile_v_3_MPORT_31_addr = 8'h23;
  assign rf_a_tile_v_3_MPORT_31_data = rf[rf_a_tile_v_3_MPORT_31_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_2_MPORT_31_en = handshaked & _GEN_1545;
  assign rf_a_tile_v_2_MPORT_31_addr = 8'h27;
  assign rf_a_tile_v_2_MPORT_31_data = rf[rf_a_tile_v_2_MPORT_31_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_1_MPORT_93_en = handshaked & _GEN_1545;
  assign rf_a_tile_v_1_MPORT_93_addr = 8'h2b;
  assign rf_a_tile_v_1_MPORT_93_data = rf[rf_a_tile_v_1_MPORT_93_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_0_MPORT_93_en = handshaked & _GEN_1545;
  assign rf_a_tile_v_0_MPORT_93_addr = 8'h2f;
  assign rf_a_tile_v_0_MPORT_93_data = rf[rf_a_tile_v_0_MPORT_93_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_3_tile_v_3_MPORT_21_en = handshaked & _GEN_1545;
  assign rf_matrix_b_3_tile_v_3_MPORT_21_addr = 8'h72;
  assign rf_matrix_b_3_tile_v_3_MPORT_21_data = rf[rf_matrix_b_3_tile_v_3_MPORT_21_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_3_tile_v_2_MPORT_21_en = handshaked & _GEN_1545;
  assign rf_matrix_b_3_tile_v_2_MPORT_21_addr = 8'h76;
  assign rf_matrix_b_3_tile_v_2_MPORT_21_data = rf[rf_matrix_b_3_tile_v_2_MPORT_21_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_3_tile_v_1_MPORT_21_en = handshaked & _GEN_1545;
  assign rf_matrix_b_3_tile_v_1_MPORT_21_addr = 8'h7a;
  assign rf_matrix_b_3_tile_v_1_MPORT_21_data = rf[rf_matrix_b_3_tile_v_1_MPORT_21_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_3_tile_v_0_MPORT_21_en = handshaked & _GEN_1545;
  assign rf_matrix_b_3_tile_v_0_MPORT_21_addr = 8'h7e;
  assign rf_matrix_b_3_tile_v_0_MPORT_21_data = rf[rf_matrix_b_3_tile_v_0_MPORT_21_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_3_tile_v_3_MPORT_21_en = handshaked & _GEN_1545;
  assign rf_matrix_c_3_tile_v_3_MPORT_21_addr = 8'ha3;
  assign rf_matrix_c_3_tile_v_3_MPORT_21_data = rf[rf_matrix_c_3_tile_v_3_MPORT_21_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_3_tile_v_2_MPORT_21_en = handshaked & _GEN_1545;
  assign rf_matrix_c_3_tile_v_2_MPORT_21_addr = 8'ha7;
  assign rf_matrix_c_3_tile_v_2_MPORT_21_data = rf[rf_matrix_c_3_tile_v_2_MPORT_21_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_3_tile_v_1_MPORT_21_en = handshaked & _GEN_1545;
  assign rf_matrix_c_3_tile_v_1_MPORT_21_addr = 8'hab;
  assign rf_matrix_c_3_tile_v_1_MPORT_21_data = rf[rf_matrix_c_3_tile_v_1_MPORT_21_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_3_tile_v_0_MPORT_21_en = handshaked & _GEN_1545;
  assign rf_matrix_c_3_tile_v_0_MPORT_21_addr = 8'haf;
  assign rf_matrix_c_3_tile_v_0_MPORT_21_data = rf[rf_matrix_c_3_tile_v_0_MPORT_21_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_1_MPORT_94_en = handshaked & _GEN_1559;
  assign rf_a_tile_v_1_MPORT_94_addr = 8'h23;
  assign rf_a_tile_v_1_MPORT_94_data = rf[rf_a_tile_v_1_MPORT_94_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_0_MPORT_94_en = handshaked & _GEN_1559;
  assign rf_a_tile_v_0_MPORT_94_addr = 8'h27;
  assign rf_a_tile_v_0_MPORT_94_data = rf[rf_a_tile_v_0_MPORT_94_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_3_tile_v_3_MPORT_22_en = handshaked & _GEN_1559;
  assign rf_matrix_b_3_tile_v_3_MPORT_22_addr = 8'h72;
  assign rf_matrix_b_3_tile_v_3_MPORT_22_data = rf[rf_matrix_b_3_tile_v_3_MPORT_22_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_3_tile_v_2_MPORT_22_en = handshaked & _GEN_1559;
  assign rf_matrix_b_3_tile_v_2_MPORT_22_addr = 8'h76;
  assign rf_matrix_b_3_tile_v_2_MPORT_22_data = rf[rf_matrix_b_3_tile_v_2_MPORT_22_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_3_tile_v_1_MPORT_22_en = handshaked & _GEN_1559;
  assign rf_matrix_b_3_tile_v_1_MPORT_22_addr = 8'h7a;
  assign rf_matrix_b_3_tile_v_1_MPORT_22_data = rf[rf_matrix_b_3_tile_v_1_MPORT_22_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_3_tile_v_0_MPORT_22_en = handshaked & _GEN_1559;
  assign rf_matrix_b_3_tile_v_0_MPORT_22_addr = 8'h7e;
  assign rf_matrix_b_3_tile_v_0_MPORT_22_data = rf[rf_matrix_b_3_tile_v_0_MPORT_22_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_3_tile_v_3_MPORT_22_en = handshaked & _GEN_1559;
  assign rf_matrix_c_3_tile_v_3_MPORT_22_addr = 8'hc6;
  assign rf_matrix_c_3_tile_v_3_MPORT_22_data = rf[rf_matrix_c_3_tile_v_3_MPORT_22_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_3_tile_v_2_MPORT_22_en = handshaked & _GEN_1559;
  assign rf_matrix_c_3_tile_v_2_MPORT_22_addr = 8'hc7;
  assign rf_matrix_c_3_tile_v_2_MPORT_22_data = rf[rf_matrix_c_3_tile_v_2_MPORT_22_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_3_tile_v_1_MPORT_22_en = handshaked & _GEN_1559;
  assign rf_matrix_c_3_tile_v_1_MPORT_22_addr = 8'hce;
  assign rf_matrix_c_3_tile_v_1_MPORT_22_data = rf[rf_matrix_c_3_tile_v_1_MPORT_22_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_3_tile_v_0_MPORT_22_en = handshaked & _GEN_1559;
  assign rf_matrix_c_3_tile_v_0_MPORT_22_addr = 8'hcf;
  assign rf_matrix_c_3_tile_v_0_MPORT_22_data = rf[rf_matrix_c_3_tile_v_0_MPORT_22_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_1_MPORT_95_en = handshaked & _GEN_1571;
  assign rf_a_tile_v_1_MPORT_95_addr = 8'h2b;
  assign rf_a_tile_v_1_MPORT_95_data = rf[rf_a_tile_v_1_MPORT_95_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_0_MPORT_95_en = handshaked & _GEN_1571;
  assign rf_a_tile_v_0_MPORT_95_addr = 8'h2f;
  assign rf_a_tile_v_0_MPORT_95_data = rf[rf_a_tile_v_0_MPORT_95_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_3_tile_v_3_MPORT_23_en = handshaked & _GEN_1571;
  assign rf_matrix_b_3_tile_v_3_MPORT_23_addr = 8'h72;
  assign rf_matrix_b_3_tile_v_3_MPORT_23_data = rf[rf_matrix_b_3_tile_v_3_MPORT_23_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_3_tile_v_2_MPORT_23_en = handshaked & _GEN_1571;
  assign rf_matrix_b_3_tile_v_2_MPORT_23_addr = 8'h76;
  assign rf_matrix_b_3_tile_v_2_MPORT_23_data = rf[rf_matrix_b_3_tile_v_2_MPORT_23_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_3_tile_v_1_MPORT_23_en = handshaked & _GEN_1571;
  assign rf_matrix_b_3_tile_v_1_MPORT_23_addr = 8'h7a;
  assign rf_matrix_b_3_tile_v_1_MPORT_23_data = rf[rf_matrix_b_3_tile_v_1_MPORT_23_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_3_tile_v_0_MPORT_23_en = handshaked & _GEN_1571;
  assign rf_matrix_b_3_tile_v_0_MPORT_23_addr = 8'h7e;
  assign rf_matrix_b_3_tile_v_0_MPORT_23_data = rf[rf_matrix_b_3_tile_v_0_MPORT_23_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_3_tile_v_3_MPORT_23_en = handshaked & _GEN_1571;
  assign rf_matrix_c_3_tile_v_3_MPORT_23_addr = 8'hd6;
  assign rf_matrix_c_3_tile_v_3_MPORT_23_data = rf[rf_matrix_c_3_tile_v_3_MPORT_23_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_3_tile_v_2_MPORT_23_en = handshaked & _GEN_1571;
  assign rf_matrix_c_3_tile_v_2_MPORT_23_addr = 8'hd7;
  assign rf_matrix_c_3_tile_v_2_MPORT_23_data = rf[rf_matrix_c_3_tile_v_2_MPORT_23_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_3_tile_v_1_MPORT_23_en = handshaked & _GEN_1571;
  assign rf_matrix_c_3_tile_v_1_MPORT_23_addr = 8'hde;
  assign rf_matrix_c_3_tile_v_1_MPORT_23_data = rf[rf_matrix_c_3_tile_v_1_MPORT_23_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_3_tile_v_0_MPORT_23_en = handshaked & _GEN_1571;
  assign rf_matrix_c_3_tile_v_0_MPORT_23_addr = 8'hdf;
  assign rf_matrix_c_3_tile_v_0_MPORT_23_data = rf[rf_matrix_c_3_tile_v_0_MPORT_23_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_1_MPORT_96_en = handshaked & _GEN_1276;
  assign rf_a_tile_v_1_MPORT_96_addr = 8'h10;
  assign rf_a_tile_v_1_MPORT_96_data = rf[rf_a_tile_v_1_MPORT_96_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_0_MPORT_96_en = handshaked & _GEN_1276;
  assign rf_a_tile_v_0_MPORT_96_addr = 8'h14;
  assign rf_a_tile_v_0_MPORT_96_data = rf[rf_a_tile_v_0_MPORT_96_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_4_tile_v_3_MPORT_en = handshaked & _GEN_1276;
  assign rf_matrix_b_4_tile_v_3_MPORT_addr = 8'h41;
  assign rf_matrix_b_4_tile_v_3_MPORT_data = rf[rf_matrix_b_4_tile_v_3_MPORT_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_4_tile_v_2_MPORT_en = handshaked & _GEN_1276;
  assign rf_matrix_b_4_tile_v_2_MPORT_addr = 8'h45;
  assign rf_matrix_b_4_tile_v_2_MPORT_data = rf[rf_matrix_b_4_tile_v_2_MPORT_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_4_tile_v_1_MPORT_en = handshaked & _GEN_1276;
  assign rf_matrix_b_4_tile_v_1_MPORT_addr = 8'h49;
  assign rf_matrix_b_4_tile_v_1_MPORT_data = rf[rf_matrix_b_4_tile_v_1_MPORT_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_4_tile_v_0_MPORT_en = handshaked & _GEN_1276;
  assign rf_matrix_b_4_tile_v_0_MPORT_addr = 8'h4d;
  assign rf_matrix_b_4_tile_v_0_MPORT_data = rf[rf_matrix_b_4_tile_v_0_MPORT_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_4_tile_v_3_MPORT_en = handshaked & _GEN_1276;
  assign rf_matrix_c_4_tile_v_3_MPORT_addr = 8'ha0;
  assign rf_matrix_c_4_tile_v_3_MPORT_data = rf[rf_matrix_c_4_tile_v_3_MPORT_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_4_tile_v_2_MPORT_en = handshaked & _GEN_1276;
  assign rf_matrix_c_4_tile_v_2_MPORT_addr = 8'ha1;
  assign rf_matrix_c_4_tile_v_2_MPORT_data = rf[rf_matrix_c_4_tile_v_2_MPORT_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_4_tile_v_1_MPORT_en = handshaked & _GEN_1276;
  assign rf_matrix_c_4_tile_v_1_MPORT_addr = 8'ha8;
  assign rf_matrix_c_4_tile_v_1_MPORT_data = rf[rf_matrix_c_4_tile_v_1_MPORT_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_4_tile_v_0_MPORT_en = handshaked & _GEN_1276;
  assign rf_matrix_c_4_tile_v_0_MPORT_addr = 8'ha9;
  assign rf_matrix_c_4_tile_v_0_MPORT_data = rf[rf_matrix_c_4_tile_v_0_MPORT_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_3_MPORT_32_en = handshaked & _GEN_1291;
  assign rf_a_tile_v_3_MPORT_32_addr = 8'h10;
  assign rf_a_tile_v_3_MPORT_32_data = rf[rf_a_tile_v_3_MPORT_32_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_2_MPORT_32_en = handshaked & _GEN_1291;
  assign rf_a_tile_v_2_MPORT_32_addr = 8'h14;
  assign rf_a_tile_v_2_MPORT_32_data = rf[rf_a_tile_v_2_MPORT_32_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_1_MPORT_97_en = handshaked & _GEN_1291;
  assign rf_a_tile_v_1_MPORT_97_addr = 8'h18;
  assign rf_a_tile_v_1_MPORT_97_data = rf[rf_a_tile_v_1_MPORT_97_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_0_MPORT_97_en = handshaked & _GEN_1291;
  assign rf_a_tile_v_0_MPORT_97_addr = 8'h1c;
  assign rf_a_tile_v_0_MPORT_97_data = rf[rf_a_tile_v_0_MPORT_97_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_4_tile_v_3_MPORT_1_en = handshaked & _GEN_1291;
  assign rf_matrix_b_4_tile_v_3_MPORT_1_addr = 8'h41;
  assign rf_matrix_b_4_tile_v_3_MPORT_1_data = rf[rf_matrix_b_4_tile_v_3_MPORT_1_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_4_tile_v_2_MPORT_1_en = handshaked & _GEN_1291;
  assign rf_matrix_b_4_tile_v_2_MPORT_1_addr = 8'h45;
  assign rf_matrix_b_4_tile_v_2_MPORT_1_data = rf[rf_matrix_b_4_tile_v_2_MPORT_1_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_4_tile_v_1_MPORT_1_en = handshaked & _GEN_1291;
  assign rf_matrix_b_4_tile_v_1_MPORT_1_addr = 8'h49;
  assign rf_matrix_b_4_tile_v_1_MPORT_1_data = rf[rf_matrix_b_4_tile_v_1_MPORT_1_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_4_tile_v_0_MPORT_1_en = handshaked & _GEN_1291;
  assign rf_matrix_b_4_tile_v_0_MPORT_1_addr = 8'h4d;
  assign rf_matrix_b_4_tile_v_0_MPORT_1_data = rf[rf_matrix_b_4_tile_v_0_MPORT_1_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_4_tile_v_3_MPORT_1_en = handshaked & _GEN_1291;
  assign rf_matrix_c_4_tile_v_3_MPORT_1_addr = 8'h90;
  assign rf_matrix_c_4_tile_v_3_MPORT_1_data = rf[rf_matrix_c_4_tile_v_3_MPORT_1_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_4_tile_v_2_MPORT_1_en = handshaked & _GEN_1291;
  assign rf_matrix_c_4_tile_v_2_MPORT_1_addr = 8'h94;
  assign rf_matrix_c_4_tile_v_2_MPORT_1_data = rf[rf_matrix_c_4_tile_v_2_MPORT_1_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_4_tile_v_1_MPORT_1_en = handshaked & _GEN_1291;
  assign rf_matrix_c_4_tile_v_1_MPORT_1_addr = 8'h98;
  assign rf_matrix_c_4_tile_v_1_MPORT_1_data = rf[rf_matrix_c_4_tile_v_1_MPORT_1_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_4_tile_v_0_MPORT_1_en = handshaked & _GEN_1291;
  assign rf_matrix_c_4_tile_v_0_MPORT_1_addr = 8'h9c;
  assign rf_matrix_c_4_tile_v_0_MPORT_1_data = rf[rf_matrix_c_4_tile_v_0_MPORT_1_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_1_MPORT_98_en = handshaked & _GEN_1305;
  assign rf_a_tile_v_1_MPORT_98_addr = 8'h18;
  assign rf_a_tile_v_1_MPORT_98_data = rf[rf_a_tile_v_1_MPORT_98_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_0_MPORT_98_en = handshaked & _GEN_1305;
  assign rf_a_tile_v_0_MPORT_98_addr = 8'h1c;
  assign rf_a_tile_v_0_MPORT_98_data = rf[rf_a_tile_v_0_MPORT_98_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_4_tile_v_3_MPORT_2_en = handshaked & _GEN_1305;
  assign rf_matrix_b_4_tile_v_3_MPORT_2_addr = 8'h41;
  assign rf_matrix_b_4_tile_v_3_MPORT_2_data = rf[rf_matrix_b_4_tile_v_3_MPORT_2_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_4_tile_v_2_MPORT_2_en = handshaked & _GEN_1305;
  assign rf_matrix_b_4_tile_v_2_MPORT_2_addr = 8'h45;
  assign rf_matrix_b_4_tile_v_2_MPORT_2_data = rf[rf_matrix_b_4_tile_v_2_MPORT_2_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_4_tile_v_1_MPORT_2_en = handshaked & _GEN_1305;
  assign rf_matrix_b_4_tile_v_1_MPORT_2_addr = 8'h49;
  assign rf_matrix_b_4_tile_v_1_MPORT_2_data = rf[rf_matrix_b_4_tile_v_1_MPORT_2_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_4_tile_v_0_MPORT_2_en = handshaked & _GEN_1305;
  assign rf_matrix_b_4_tile_v_0_MPORT_2_addr = 8'h4d;
  assign rf_matrix_b_4_tile_v_0_MPORT_2_data = rf[rf_matrix_b_4_tile_v_0_MPORT_2_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_4_tile_v_3_MPORT_2_en = handshaked & _GEN_1305;
  assign rf_matrix_c_4_tile_v_3_MPORT_2_addr = 8'hb0;
  assign rf_matrix_c_4_tile_v_3_MPORT_2_data = rf[rf_matrix_c_4_tile_v_3_MPORT_2_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_4_tile_v_2_MPORT_2_en = handshaked & _GEN_1305;
  assign rf_matrix_c_4_tile_v_2_MPORT_2_addr = 8'hb1;
  assign rf_matrix_c_4_tile_v_2_MPORT_2_data = rf[rf_matrix_c_4_tile_v_2_MPORT_2_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_4_tile_v_1_MPORT_2_en = handshaked & _GEN_1305;
  assign rf_matrix_c_4_tile_v_1_MPORT_2_addr = 8'hb8;
  assign rf_matrix_c_4_tile_v_1_MPORT_2_data = rf[rf_matrix_c_4_tile_v_1_MPORT_2_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_4_tile_v_0_MPORT_2_en = handshaked & _GEN_1305;
  assign rf_matrix_c_4_tile_v_0_MPORT_2_addr = 8'hb9;
  assign rf_matrix_c_4_tile_v_0_MPORT_2_data = rf[rf_matrix_c_4_tile_v_0_MPORT_2_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_3_MPORT_33_en = handshaked & _GEN_1317;
  assign rf_a_tile_v_3_MPORT_33_addr = 8'h10;
  assign rf_a_tile_v_3_MPORT_33_data = rf[rf_a_tile_v_3_MPORT_33_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_2_MPORT_33_en = handshaked & _GEN_1317;
  assign rf_a_tile_v_2_MPORT_33_addr = 8'h14;
  assign rf_a_tile_v_2_MPORT_33_data = rf[rf_a_tile_v_2_MPORT_33_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_1_MPORT_99_en = handshaked & _GEN_1317;
  assign rf_a_tile_v_1_MPORT_99_addr = 8'h18;
  assign rf_a_tile_v_1_MPORT_99_data = rf[rf_a_tile_v_1_MPORT_99_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_0_MPORT_99_en = handshaked & _GEN_1317;
  assign rf_a_tile_v_0_MPORT_99_addr = 8'h1c;
  assign rf_a_tile_v_0_MPORT_99_data = rf[rf_a_tile_v_0_MPORT_99_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_4_tile_v_3_MPORT_3_en = handshaked & _GEN_1317;
  assign rf_matrix_b_4_tile_v_3_MPORT_3_addr = 8'h41;
  assign rf_matrix_b_4_tile_v_3_MPORT_3_data = rf[rf_matrix_b_4_tile_v_3_MPORT_3_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_4_tile_v_2_MPORT_3_en = handshaked & _GEN_1317;
  assign rf_matrix_b_4_tile_v_2_MPORT_3_addr = 8'h45;
  assign rf_matrix_b_4_tile_v_2_MPORT_3_data = rf[rf_matrix_b_4_tile_v_2_MPORT_3_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_4_tile_v_1_MPORT_3_en = handshaked & _GEN_1317;
  assign rf_matrix_b_4_tile_v_1_MPORT_3_addr = 8'h49;
  assign rf_matrix_b_4_tile_v_1_MPORT_3_data = rf[rf_matrix_b_4_tile_v_1_MPORT_3_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_4_tile_v_0_MPORT_3_en = handshaked & _GEN_1317;
  assign rf_matrix_b_4_tile_v_0_MPORT_3_addr = 8'h4d;
  assign rf_matrix_b_4_tile_v_0_MPORT_3_data = rf[rf_matrix_b_4_tile_v_0_MPORT_3_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_4_tile_v_3_MPORT_3_en = handshaked & _GEN_1317;
  assign rf_matrix_c_4_tile_v_3_MPORT_3_addr = 8'h91;
  assign rf_matrix_c_4_tile_v_3_MPORT_3_data = rf[rf_matrix_c_4_tile_v_3_MPORT_3_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_4_tile_v_2_MPORT_3_en = handshaked & _GEN_1317;
  assign rf_matrix_c_4_tile_v_2_MPORT_3_addr = 8'h95;
  assign rf_matrix_c_4_tile_v_2_MPORT_3_data = rf[rf_matrix_c_4_tile_v_2_MPORT_3_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_4_tile_v_1_MPORT_3_en = handshaked & _GEN_1317;
  assign rf_matrix_c_4_tile_v_1_MPORT_3_addr = 8'h99;
  assign rf_matrix_c_4_tile_v_1_MPORT_3_data = rf[rf_matrix_c_4_tile_v_1_MPORT_3_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_4_tile_v_0_MPORT_3_en = handshaked & _GEN_1317;
  assign rf_matrix_c_4_tile_v_0_MPORT_3_addr = 8'h9d;
  assign rf_matrix_c_4_tile_v_0_MPORT_3_data = rf[rf_matrix_c_4_tile_v_0_MPORT_3_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_1_MPORT_100_en = handshaked & _GEN_1331;
  assign rf_a_tile_v_1_MPORT_100_addr = 8'h10;
  assign rf_a_tile_v_1_MPORT_100_data = rf[rf_a_tile_v_1_MPORT_100_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_0_MPORT_100_en = handshaked & _GEN_1331;
  assign rf_a_tile_v_0_MPORT_100_addr = 8'h14;
  assign rf_a_tile_v_0_MPORT_100_data = rf[rf_a_tile_v_0_MPORT_100_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_4_tile_v_3_MPORT_4_en = handshaked & _GEN_1331;
  assign rf_matrix_b_4_tile_v_3_MPORT_4_addr = 8'h41;
  assign rf_matrix_b_4_tile_v_3_MPORT_4_data = rf[rf_matrix_b_4_tile_v_3_MPORT_4_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_4_tile_v_2_MPORT_4_en = handshaked & _GEN_1331;
  assign rf_matrix_b_4_tile_v_2_MPORT_4_addr = 8'h45;
  assign rf_matrix_b_4_tile_v_2_MPORT_4_data = rf[rf_matrix_b_4_tile_v_2_MPORT_4_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_4_tile_v_1_MPORT_4_en = handshaked & _GEN_1331;
  assign rf_matrix_b_4_tile_v_1_MPORT_4_addr = 8'h49;
  assign rf_matrix_b_4_tile_v_1_MPORT_4_data = rf[rf_matrix_b_4_tile_v_1_MPORT_4_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_4_tile_v_0_MPORT_4_en = handshaked & _GEN_1331;
  assign rf_matrix_b_4_tile_v_0_MPORT_4_addr = 8'h4d;
  assign rf_matrix_b_4_tile_v_0_MPORT_4_data = rf[rf_matrix_b_4_tile_v_0_MPORT_4_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_4_tile_v_3_MPORT_4_en = handshaked & _GEN_1331;
  assign rf_matrix_c_4_tile_v_3_MPORT_4_addr = 8'ha2;
  assign rf_matrix_c_4_tile_v_3_MPORT_4_data = rf[rf_matrix_c_4_tile_v_3_MPORT_4_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_4_tile_v_2_MPORT_4_en = handshaked & _GEN_1331;
  assign rf_matrix_c_4_tile_v_2_MPORT_4_addr = 8'ha3;
  assign rf_matrix_c_4_tile_v_2_MPORT_4_data = rf[rf_matrix_c_4_tile_v_2_MPORT_4_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_4_tile_v_1_MPORT_4_en = handshaked & _GEN_1331;
  assign rf_matrix_c_4_tile_v_1_MPORT_4_addr = 8'haa;
  assign rf_matrix_c_4_tile_v_1_MPORT_4_data = rf[rf_matrix_c_4_tile_v_1_MPORT_4_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_4_tile_v_0_MPORT_4_en = handshaked & _GEN_1331;
  assign rf_matrix_c_4_tile_v_0_MPORT_4_addr = 8'hab;
  assign rf_matrix_c_4_tile_v_0_MPORT_4_data = rf[rf_matrix_c_4_tile_v_0_MPORT_4_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_1_MPORT_101_en = handshaked & _GEN_1343;
  assign rf_a_tile_v_1_MPORT_101_addr = 8'h18;
  assign rf_a_tile_v_1_MPORT_101_data = rf[rf_a_tile_v_1_MPORT_101_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_0_MPORT_101_en = handshaked & _GEN_1343;
  assign rf_a_tile_v_0_MPORT_101_addr = 8'h1c;
  assign rf_a_tile_v_0_MPORT_101_data = rf[rf_a_tile_v_0_MPORT_101_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_4_tile_v_3_MPORT_5_en = handshaked & _GEN_1343;
  assign rf_matrix_b_4_tile_v_3_MPORT_5_addr = 8'h41;
  assign rf_matrix_b_4_tile_v_3_MPORT_5_data = rf[rf_matrix_b_4_tile_v_3_MPORT_5_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_4_tile_v_2_MPORT_5_en = handshaked & _GEN_1343;
  assign rf_matrix_b_4_tile_v_2_MPORT_5_addr = 8'h45;
  assign rf_matrix_b_4_tile_v_2_MPORT_5_data = rf[rf_matrix_b_4_tile_v_2_MPORT_5_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_4_tile_v_1_MPORT_5_en = handshaked & _GEN_1343;
  assign rf_matrix_b_4_tile_v_1_MPORT_5_addr = 8'h49;
  assign rf_matrix_b_4_tile_v_1_MPORT_5_data = rf[rf_matrix_b_4_tile_v_1_MPORT_5_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_4_tile_v_0_MPORT_5_en = handshaked & _GEN_1343;
  assign rf_matrix_b_4_tile_v_0_MPORT_5_addr = 8'h4d;
  assign rf_matrix_b_4_tile_v_0_MPORT_5_data = rf[rf_matrix_b_4_tile_v_0_MPORT_5_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_4_tile_v_3_MPORT_5_en = handshaked & _GEN_1343;
  assign rf_matrix_c_4_tile_v_3_MPORT_5_addr = 8'hb2;
  assign rf_matrix_c_4_tile_v_3_MPORT_5_data = rf[rf_matrix_c_4_tile_v_3_MPORT_5_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_4_tile_v_2_MPORT_5_en = handshaked & _GEN_1343;
  assign rf_matrix_c_4_tile_v_2_MPORT_5_addr = 8'hb3;
  assign rf_matrix_c_4_tile_v_2_MPORT_5_data = rf[rf_matrix_c_4_tile_v_2_MPORT_5_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_4_tile_v_1_MPORT_5_en = handshaked & _GEN_1343;
  assign rf_matrix_c_4_tile_v_1_MPORT_5_addr = 8'hba;
  assign rf_matrix_c_4_tile_v_1_MPORT_5_data = rf[rf_matrix_c_4_tile_v_1_MPORT_5_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_4_tile_v_0_MPORT_5_en = handshaked & _GEN_1343;
  assign rf_matrix_c_4_tile_v_0_MPORT_5_addr = 8'hbb;
  assign rf_matrix_c_4_tile_v_0_MPORT_5_data = rf[rf_matrix_c_4_tile_v_0_MPORT_5_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_1_MPORT_102_en = handshaked & _GEN_1355;
  assign rf_a_tile_v_1_MPORT_102_addr = 8'h11;
  assign rf_a_tile_v_1_MPORT_102_data = rf[rf_a_tile_v_1_MPORT_102_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_0_MPORT_102_en = handshaked & _GEN_1355;
  assign rf_a_tile_v_0_MPORT_102_addr = 8'h15;
  assign rf_a_tile_v_0_MPORT_102_data = rf[rf_a_tile_v_0_MPORT_102_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_4_tile_v_3_MPORT_6_en = handshaked & _GEN_1355;
  assign rf_matrix_b_4_tile_v_3_MPORT_6_addr = 8'h51;
  assign rf_matrix_b_4_tile_v_3_MPORT_6_data = rf[rf_matrix_b_4_tile_v_3_MPORT_6_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_4_tile_v_2_MPORT_6_en = handshaked & _GEN_1355;
  assign rf_matrix_b_4_tile_v_2_MPORT_6_addr = 8'h55;
  assign rf_matrix_b_4_tile_v_2_MPORT_6_data = rf[rf_matrix_b_4_tile_v_2_MPORT_6_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_4_tile_v_1_MPORT_6_en = handshaked & _GEN_1355;
  assign rf_matrix_b_4_tile_v_1_MPORT_6_addr = 8'h59;
  assign rf_matrix_b_4_tile_v_1_MPORT_6_data = rf[rf_matrix_b_4_tile_v_1_MPORT_6_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_4_tile_v_0_MPORT_6_en = handshaked & _GEN_1355;
  assign rf_matrix_b_4_tile_v_0_MPORT_6_addr = 8'h5d;
  assign rf_matrix_b_4_tile_v_0_MPORT_6_data = rf[rf_matrix_b_4_tile_v_0_MPORT_6_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_4_tile_v_3_MPORT_6_en = handshaked & _GEN_1355;
  assign rf_matrix_c_4_tile_v_3_MPORT_6_addr = 8'ha0;
  assign rf_matrix_c_4_tile_v_3_MPORT_6_data = rf[rf_matrix_c_4_tile_v_3_MPORT_6_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_4_tile_v_2_MPORT_6_en = handshaked & _GEN_1355;
  assign rf_matrix_c_4_tile_v_2_MPORT_6_addr = 8'ha1;
  assign rf_matrix_c_4_tile_v_2_MPORT_6_data = rf[rf_matrix_c_4_tile_v_2_MPORT_6_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_4_tile_v_1_MPORT_6_en = handshaked & _GEN_1355;
  assign rf_matrix_c_4_tile_v_1_MPORT_6_addr = 8'ha8;
  assign rf_matrix_c_4_tile_v_1_MPORT_6_data = rf[rf_matrix_c_4_tile_v_1_MPORT_6_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_4_tile_v_0_MPORT_6_en = handshaked & _GEN_1355;
  assign rf_matrix_c_4_tile_v_0_MPORT_6_addr = 8'ha9;
  assign rf_matrix_c_4_tile_v_0_MPORT_6_data = rf[rf_matrix_c_4_tile_v_0_MPORT_6_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_3_MPORT_34_en = handshaked & _GEN_1367;
  assign rf_a_tile_v_3_MPORT_34_addr = 8'h11;
  assign rf_a_tile_v_3_MPORT_34_data = rf[rf_a_tile_v_3_MPORT_34_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_2_MPORT_34_en = handshaked & _GEN_1367;
  assign rf_a_tile_v_2_MPORT_34_addr = 8'h15;
  assign rf_a_tile_v_2_MPORT_34_data = rf[rf_a_tile_v_2_MPORT_34_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_1_MPORT_103_en = handshaked & _GEN_1367;
  assign rf_a_tile_v_1_MPORT_103_addr = 8'h19;
  assign rf_a_tile_v_1_MPORT_103_data = rf[rf_a_tile_v_1_MPORT_103_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_0_MPORT_103_en = handshaked & _GEN_1367;
  assign rf_a_tile_v_0_MPORT_103_addr = 8'h1d;
  assign rf_a_tile_v_0_MPORT_103_data = rf[rf_a_tile_v_0_MPORT_103_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_4_tile_v_3_MPORT_7_en = handshaked & _GEN_1367;
  assign rf_matrix_b_4_tile_v_3_MPORT_7_addr = 8'h51;
  assign rf_matrix_b_4_tile_v_3_MPORT_7_data = rf[rf_matrix_b_4_tile_v_3_MPORT_7_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_4_tile_v_2_MPORT_7_en = handshaked & _GEN_1367;
  assign rf_matrix_b_4_tile_v_2_MPORT_7_addr = 8'h55;
  assign rf_matrix_b_4_tile_v_2_MPORT_7_data = rf[rf_matrix_b_4_tile_v_2_MPORT_7_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_4_tile_v_1_MPORT_7_en = handshaked & _GEN_1367;
  assign rf_matrix_b_4_tile_v_1_MPORT_7_addr = 8'h59;
  assign rf_matrix_b_4_tile_v_1_MPORT_7_data = rf[rf_matrix_b_4_tile_v_1_MPORT_7_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_4_tile_v_0_MPORT_7_en = handshaked & _GEN_1367;
  assign rf_matrix_b_4_tile_v_0_MPORT_7_addr = 8'h5d;
  assign rf_matrix_b_4_tile_v_0_MPORT_7_data = rf[rf_matrix_b_4_tile_v_0_MPORT_7_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_4_tile_v_3_MPORT_7_en = handshaked & _GEN_1367;
  assign rf_matrix_c_4_tile_v_3_MPORT_7_addr = 8'h90;
  assign rf_matrix_c_4_tile_v_3_MPORT_7_data = rf[rf_matrix_c_4_tile_v_3_MPORT_7_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_4_tile_v_2_MPORT_7_en = handshaked & _GEN_1367;
  assign rf_matrix_c_4_tile_v_2_MPORT_7_addr = 8'h94;
  assign rf_matrix_c_4_tile_v_2_MPORT_7_data = rf[rf_matrix_c_4_tile_v_2_MPORT_7_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_4_tile_v_1_MPORT_7_en = handshaked & _GEN_1367;
  assign rf_matrix_c_4_tile_v_1_MPORT_7_addr = 8'h98;
  assign rf_matrix_c_4_tile_v_1_MPORT_7_data = rf[rf_matrix_c_4_tile_v_1_MPORT_7_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_4_tile_v_0_MPORT_7_en = handshaked & _GEN_1367;
  assign rf_matrix_c_4_tile_v_0_MPORT_7_addr = 8'h9c;
  assign rf_matrix_c_4_tile_v_0_MPORT_7_data = rf[rf_matrix_c_4_tile_v_0_MPORT_7_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_1_MPORT_104_en = handshaked & _GEN_1381;
  assign rf_a_tile_v_1_MPORT_104_addr = 8'h19;
  assign rf_a_tile_v_1_MPORT_104_data = rf[rf_a_tile_v_1_MPORT_104_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_0_MPORT_104_en = handshaked & _GEN_1381;
  assign rf_a_tile_v_0_MPORT_104_addr = 8'h1d;
  assign rf_a_tile_v_0_MPORT_104_data = rf[rf_a_tile_v_0_MPORT_104_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_4_tile_v_3_MPORT_8_en = handshaked & _GEN_1381;
  assign rf_matrix_b_4_tile_v_3_MPORT_8_addr = 8'h51;
  assign rf_matrix_b_4_tile_v_3_MPORT_8_data = rf[rf_matrix_b_4_tile_v_3_MPORT_8_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_4_tile_v_2_MPORT_8_en = handshaked & _GEN_1381;
  assign rf_matrix_b_4_tile_v_2_MPORT_8_addr = 8'h55;
  assign rf_matrix_b_4_tile_v_2_MPORT_8_data = rf[rf_matrix_b_4_tile_v_2_MPORT_8_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_4_tile_v_1_MPORT_8_en = handshaked & _GEN_1381;
  assign rf_matrix_b_4_tile_v_1_MPORT_8_addr = 8'h59;
  assign rf_matrix_b_4_tile_v_1_MPORT_8_data = rf[rf_matrix_b_4_tile_v_1_MPORT_8_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_4_tile_v_0_MPORT_8_en = handshaked & _GEN_1381;
  assign rf_matrix_b_4_tile_v_0_MPORT_8_addr = 8'h5d;
  assign rf_matrix_b_4_tile_v_0_MPORT_8_data = rf[rf_matrix_b_4_tile_v_0_MPORT_8_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_4_tile_v_3_MPORT_8_en = handshaked & _GEN_1381;
  assign rf_matrix_c_4_tile_v_3_MPORT_8_addr = 8'hb0;
  assign rf_matrix_c_4_tile_v_3_MPORT_8_data = rf[rf_matrix_c_4_tile_v_3_MPORT_8_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_4_tile_v_2_MPORT_8_en = handshaked & _GEN_1381;
  assign rf_matrix_c_4_tile_v_2_MPORT_8_addr = 8'hb1;
  assign rf_matrix_c_4_tile_v_2_MPORT_8_data = rf[rf_matrix_c_4_tile_v_2_MPORT_8_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_4_tile_v_1_MPORT_8_en = handshaked & _GEN_1381;
  assign rf_matrix_c_4_tile_v_1_MPORT_8_addr = 8'hb8;
  assign rf_matrix_c_4_tile_v_1_MPORT_8_data = rf[rf_matrix_c_4_tile_v_1_MPORT_8_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_4_tile_v_0_MPORT_8_en = handshaked & _GEN_1381;
  assign rf_matrix_c_4_tile_v_0_MPORT_8_addr = 8'hb9;
  assign rf_matrix_c_4_tile_v_0_MPORT_8_data = rf[rf_matrix_c_4_tile_v_0_MPORT_8_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_3_MPORT_35_en = handshaked & _GEN_1393;
  assign rf_a_tile_v_3_MPORT_35_addr = 8'h11;
  assign rf_a_tile_v_3_MPORT_35_data = rf[rf_a_tile_v_3_MPORT_35_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_2_MPORT_35_en = handshaked & _GEN_1393;
  assign rf_a_tile_v_2_MPORT_35_addr = 8'h15;
  assign rf_a_tile_v_2_MPORT_35_data = rf[rf_a_tile_v_2_MPORT_35_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_1_MPORT_105_en = handshaked & _GEN_1393;
  assign rf_a_tile_v_1_MPORT_105_addr = 8'h19;
  assign rf_a_tile_v_1_MPORT_105_data = rf[rf_a_tile_v_1_MPORT_105_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_0_MPORT_105_en = handshaked & _GEN_1393;
  assign rf_a_tile_v_0_MPORT_105_addr = 8'h1d;
  assign rf_a_tile_v_0_MPORT_105_data = rf[rf_a_tile_v_0_MPORT_105_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_4_tile_v_3_MPORT_9_en = handshaked & _GEN_1393;
  assign rf_matrix_b_4_tile_v_3_MPORT_9_addr = 8'h51;
  assign rf_matrix_b_4_tile_v_3_MPORT_9_data = rf[rf_matrix_b_4_tile_v_3_MPORT_9_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_4_tile_v_2_MPORT_9_en = handshaked & _GEN_1393;
  assign rf_matrix_b_4_tile_v_2_MPORT_9_addr = 8'h55;
  assign rf_matrix_b_4_tile_v_2_MPORT_9_data = rf[rf_matrix_b_4_tile_v_2_MPORT_9_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_4_tile_v_1_MPORT_9_en = handshaked & _GEN_1393;
  assign rf_matrix_b_4_tile_v_1_MPORT_9_addr = 8'h59;
  assign rf_matrix_b_4_tile_v_1_MPORT_9_data = rf[rf_matrix_b_4_tile_v_1_MPORT_9_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_4_tile_v_0_MPORT_9_en = handshaked & _GEN_1393;
  assign rf_matrix_b_4_tile_v_0_MPORT_9_addr = 8'h5d;
  assign rf_matrix_b_4_tile_v_0_MPORT_9_data = rf[rf_matrix_b_4_tile_v_0_MPORT_9_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_4_tile_v_3_MPORT_9_en = handshaked & _GEN_1393;
  assign rf_matrix_c_4_tile_v_3_MPORT_9_addr = 8'h91;
  assign rf_matrix_c_4_tile_v_3_MPORT_9_data = rf[rf_matrix_c_4_tile_v_3_MPORT_9_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_4_tile_v_2_MPORT_9_en = handshaked & _GEN_1393;
  assign rf_matrix_c_4_tile_v_2_MPORT_9_addr = 8'h95;
  assign rf_matrix_c_4_tile_v_2_MPORT_9_data = rf[rf_matrix_c_4_tile_v_2_MPORT_9_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_4_tile_v_1_MPORT_9_en = handshaked & _GEN_1393;
  assign rf_matrix_c_4_tile_v_1_MPORT_9_addr = 8'h99;
  assign rf_matrix_c_4_tile_v_1_MPORT_9_data = rf[rf_matrix_c_4_tile_v_1_MPORT_9_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_4_tile_v_0_MPORT_9_en = handshaked & _GEN_1393;
  assign rf_matrix_c_4_tile_v_0_MPORT_9_addr = 8'h9d;
  assign rf_matrix_c_4_tile_v_0_MPORT_9_data = rf[rf_matrix_c_4_tile_v_0_MPORT_9_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_1_MPORT_106_en = handshaked & _GEN_1407;
  assign rf_a_tile_v_1_MPORT_106_addr = 8'h11;
  assign rf_a_tile_v_1_MPORT_106_data = rf[rf_a_tile_v_1_MPORT_106_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_0_MPORT_106_en = handshaked & _GEN_1407;
  assign rf_a_tile_v_0_MPORT_106_addr = 8'h15;
  assign rf_a_tile_v_0_MPORT_106_data = rf[rf_a_tile_v_0_MPORT_106_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_4_tile_v_3_MPORT_10_en = handshaked & _GEN_1407;
  assign rf_matrix_b_4_tile_v_3_MPORT_10_addr = 8'h51;
  assign rf_matrix_b_4_tile_v_3_MPORT_10_data = rf[rf_matrix_b_4_tile_v_3_MPORT_10_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_4_tile_v_2_MPORT_10_en = handshaked & _GEN_1407;
  assign rf_matrix_b_4_tile_v_2_MPORT_10_addr = 8'h55;
  assign rf_matrix_b_4_tile_v_2_MPORT_10_data = rf[rf_matrix_b_4_tile_v_2_MPORT_10_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_4_tile_v_1_MPORT_10_en = handshaked & _GEN_1407;
  assign rf_matrix_b_4_tile_v_1_MPORT_10_addr = 8'h59;
  assign rf_matrix_b_4_tile_v_1_MPORT_10_data = rf[rf_matrix_b_4_tile_v_1_MPORT_10_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_4_tile_v_0_MPORT_10_en = handshaked & _GEN_1407;
  assign rf_matrix_b_4_tile_v_0_MPORT_10_addr = 8'h5d;
  assign rf_matrix_b_4_tile_v_0_MPORT_10_data = rf[rf_matrix_b_4_tile_v_0_MPORT_10_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_4_tile_v_3_MPORT_10_en = handshaked & _GEN_1407;
  assign rf_matrix_c_4_tile_v_3_MPORT_10_addr = 8'ha2;
  assign rf_matrix_c_4_tile_v_3_MPORT_10_data = rf[rf_matrix_c_4_tile_v_3_MPORT_10_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_4_tile_v_2_MPORT_10_en = handshaked & _GEN_1407;
  assign rf_matrix_c_4_tile_v_2_MPORT_10_addr = 8'ha3;
  assign rf_matrix_c_4_tile_v_2_MPORT_10_data = rf[rf_matrix_c_4_tile_v_2_MPORT_10_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_4_tile_v_1_MPORT_10_en = handshaked & _GEN_1407;
  assign rf_matrix_c_4_tile_v_1_MPORT_10_addr = 8'haa;
  assign rf_matrix_c_4_tile_v_1_MPORT_10_data = rf[rf_matrix_c_4_tile_v_1_MPORT_10_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_4_tile_v_0_MPORT_10_en = handshaked & _GEN_1407;
  assign rf_matrix_c_4_tile_v_0_MPORT_10_addr = 8'hab;
  assign rf_matrix_c_4_tile_v_0_MPORT_10_data = rf[rf_matrix_c_4_tile_v_0_MPORT_10_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_1_MPORT_107_en = handshaked & _GEN_1419;
  assign rf_a_tile_v_1_MPORT_107_addr = 8'h19;
  assign rf_a_tile_v_1_MPORT_107_data = rf[rf_a_tile_v_1_MPORT_107_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_0_MPORT_107_en = handshaked & _GEN_1419;
  assign rf_a_tile_v_0_MPORT_107_addr = 8'h1d;
  assign rf_a_tile_v_0_MPORT_107_data = rf[rf_a_tile_v_0_MPORT_107_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_4_tile_v_3_MPORT_11_en = handshaked & _GEN_1419;
  assign rf_matrix_b_4_tile_v_3_MPORT_11_addr = 8'h51;
  assign rf_matrix_b_4_tile_v_3_MPORT_11_data = rf[rf_matrix_b_4_tile_v_3_MPORT_11_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_4_tile_v_2_MPORT_11_en = handshaked & _GEN_1419;
  assign rf_matrix_b_4_tile_v_2_MPORT_11_addr = 8'h55;
  assign rf_matrix_b_4_tile_v_2_MPORT_11_data = rf[rf_matrix_b_4_tile_v_2_MPORT_11_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_4_tile_v_1_MPORT_11_en = handshaked & _GEN_1419;
  assign rf_matrix_b_4_tile_v_1_MPORT_11_addr = 8'h59;
  assign rf_matrix_b_4_tile_v_1_MPORT_11_data = rf[rf_matrix_b_4_tile_v_1_MPORT_11_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_4_tile_v_0_MPORT_11_en = handshaked & _GEN_1419;
  assign rf_matrix_b_4_tile_v_0_MPORT_11_addr = 8'h5d;
  assign rf_matrix_b_4_tile_v_0_MPORT_11_data = rf[rf_matrix_b_4_tile_v_0_MPORT_11_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_4_tile_v_3_MPORT_11_en = handshaked & _GEN_1419;
  assign rf_matrix_c_4_tile_v_3_MPORT_11_addr = 8'hb2;
  assign rf_matrix_c_4_tile_v_3_MPORT_11_data = rf[rf_matrix_c_4_tile_v_3_MPORT_11_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_4_tile_v_2_MPORT_11_en = handshaked & _GEN_1419;
  assign rf_matrix_c_4_tile_v_2_MPORT_11_addr = 8'hb3;
  assign rf_matrix_c_4_tile_v_2_MPORT_11_data = rf[rf_matrix_c_4_tile_v_2_MPORT_11_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_4_tile_v_1_MPORT_11_en = handshaked & _GEN_1419;
  assign rf_matrix_c_4_tile_v_1_MPORT_11_addr = 8'hba;
  assign rf_matrix_c_4_tile_v_1_MPORT_11_data = rf[rf_matrix_c_4_tile_v_1_MPORT_11_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_4_tile_v_0_MPORT_11_en = handshaked & _GEN_1419;
  assign rf_matrix_c_4_tile_v_0_MPORT_11_addr = 8'hbb;
  assign rf_matrix_c_4_tile_v_0_MPORT_11_data = rf[rf_matrix_c_4_tile_v_0_MPORT_11_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_1_MPORT_108_en = handshaked & _GEN_1431;
  assign rf_a_tile_v_1_MPORT_108_addr = 8'h12;
  assign rf_a_tile_v_1_MPORT_108_data = rf[rf_a_tile_v_1_MPORT_108_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_0_MPORT_108_en = handshaked & _GEN_1431;
  assign rf_a_tile_v_0_MPORT_108_addr = 8'h16;
  assign rf_a_tile_v_0_MPORT_108_data = rf[rf_a_tile_v_0_MPORT_108_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_4_tile_v_3_MPORT_12_en = handshaked & _GEN_1431;
  assign rf_matrix_b_4_tile_v_3_MPORT_12_addr = 8'h61;
  assign rf_matrix_b_4_tile_v_3_MPORT_12_data = rf[rf_matrix_b_4_tile_v_3_MPORT_12_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_4_tile_v_2_MPORT_12_en = handshaked & _GEN_1431;
  assign rf_matrix_b_4_tile_v_2_MPORT_12_addr = 8'h65;
  assign rf_matrix_b_4_tile_v_2_MPORT_12_data = rf[rf_matrix_b_4_tile_v_2_MPORT_12_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_4_tile_v_1_MPORT_12_en = handshaked & _GEN_1431;
  assign rf_matrix_b_4_tile_v_1_MPORT_12_addr = 8'h69;
  assign rf_matrix_b_4_tile_v_1_MPORT_12_data = rf[rf_matrix_b_4_tile_v_1_MPORT_12_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_4_tile_v_0_MPORT_12_en = handshaked & _GEN_1431;
  assign rf_matrix_b_4_tile_v_0_MPORT_12_addr = 8'h6d;
  assign rf_matrix_b_4_tile_v_0_MPORT_12_data = rf[rf_matrix_b_4_tile_v_0_MPORT_12_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_4_tile_v_3_MPORT_12_en = handshaked & _GEN_1431;
  assign rf_matrix_c_4_tile_v_3_MPORT_12_addr = 8'ha0;
  assign rf_matrix_c_4_tile_v_3_MPORT_12_data = rf[rf_matrix_c_4_tile_v_3_MPORT_12_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_4_tile_v_2_MPORT_12_en = handshaked & _GEN_1431;
  assign rf_matrix_c_4_tile_v_2_MPORT_12_addr = 8'ha1;
  assign rf_matrix_c_4_tile_v_2_MPORT_12_data = rf[rf_matrix_c_4_tile_v_2_MPORT_12_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_4_tile_v_1_MPORT_12_en = handshaked & _GEN_1431;
  assign rf_matrix_c_4_tile_v_1_MPORT_12_addr = 8'ha8;
  assign rf_matrix_c_4_tile_v_1_MPORT_12_data = rf[rf_matrix_c_4_tile_v_1_MPORT_12_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_4_tile_v_0_MPORT_12_en = handshaked & _GEN_1431;
  assign rf_matrix_c_4_tile_v_0_MPORT_12_addr = 8'ha9;
  assign rf_matrix_c_4_tile_v_0_MPORT_12_data = rf[rf_matrix_c_4_tile_v_0_MPORT_12_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_3_MPORT_36_en = handshaked & _GEN_1443;
  assign rf_a_tile_v_3_MPORT_36_addr = 8'h12;
  assign rf_a_tile_v_3_MPORT_36_data = rf[rf_a_tile_v_3_MPORT_36_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_2_MPORT_36_en = handshaked & _GEN_1443;
  assign rf_a_tile_v_2_MPORT_36_addr = 8'h16;
  assign rf_a_tile_v_2_MPORT_36_data = rf[rf_a_tile_v_2_MPORT_36_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_1_MPORT_109_en = handshaked & _GEN_1443;
  assign rf_a_tile_v_1_MPORT_109_addr = 8'h1a;
  assign rf_a_tile_v_1_MPORT_109_data = rf[rf_a_tile_v_1_MPORT_109_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_0_MPORT_109_en = handshaked & _GEN_1443;
  assign rf_a_tile_v_0_MPORT_109_addr = 8'h1e;
  assign rf_a_tile_v_0_MPORT_109_data = rf[rf_a_tile_v_0_MPORT_109_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_4_tile_v_3_MPORT_13_en = handshaked & _GEN_1443;
  assign rf_matrix_b_4_tile_v_3_MPORT_13_addr = 8'h61;
  assign rf_matrix_b_4_tile_v_3_MPORT_13_data = rf[rf_matrix_b_4_tile_v_3_MPORT_13_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_4_tile_v_2_MPORT_13_en = handshaked & _GEN_1443;
  assign rf_matrix_b_4_tile_v_2_MPORT_13_addr = 8'h65;
  assign rf_matrix_b_4_tile_v_2_MPORT_13_data = rf[rf_matrix_b_4_tile_v_2_MPORT_13_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_4_tile_v_1_MPORT_13_en = handshaked & _GEN_1443;
  assign rf_matrix_b_4_tile_v_1_MPORT_13_addr = 8'h69;
  assign rf_matrix_b_4_tile_v_1_MPORT_13_data = rf[rf_matrix_b_4_tile_v_1_MPORT_13_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_4_tile_v_0_MPORT_13_en = handshaked & _GEN_1443;
  assign rf_matrix_b_4_tile_v_0_MPORT_13_addr = 8'h6d;
  assign rf_matrix_b_4_tile_v_0_MPORT_13_data = rf[rf_matrix_b_4_tile_v_0_MPORT_13_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_4_tile_v_3_MPORT_13_en = handshaked & _GEN_1443;
  assign rf_matrix_c_4_tile_v_3_MPORT_13_addr = 8'h90;
  assign rf_matrix_c_4_tile_v_3_MPORT_13_data = rf[rf_matrix_c_4_tile_v_3_MPORT_13_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_4_tile_v_2_MPORT_13_en = handshaked & _GEN_1443;
  assign rf_matrix_c_4_tile_v_2_MPORT_13_addr = 8'h94;
  assign rf_matrix_c_4_tile_v_2_MPORT_13_data = rf[rf_matrix_c_4_tile_v_2_MPORT_13_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_4_tile_v_1_MPORT_13_en = handshaked & _GEN_1443;
  assign rf_matrix_c_4_tile_v_1_MPORT_13_addr = 8'h98;
  assign rf_matrix_c_4_tile_v_1_MPORT_13_data = rf[rf_matrix_c_4_tile_v_1_MPORT_13_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_4_tile_v_0_MPORT_13_en = handshaked & _GEN_1443;
  assign rf_matrix_c_4_tile_v_0_MPORT_13_addr = 8'h9c;
  assign rf_matrix_c_4_tile_v_0_MPORT_13_data = rf[rf_matrix_c_4_tile_v_0_MPORT_13_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_1_MPORT_110_en = handshaked & _GEN_1457;
  assign rf_a_tile_v_1_MPORT_110_addr = 8'h1a;
  assign rf_a_tile_v_1_MPORT_110_data = rf[rf_a_tile_v_1_MPORT_110_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_0_MPORT_110_en = handshaked & _GEN_1457;
  assign rf_a_tile_v_0_MPORT_110_addr = 8'h1e;
  assign rf_a_tile_v_0_MPORT_110_data = rf[rf_a_tile_v_0_MPORT_110_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_4_tile_v_3_MPORT_14_en = handshaked & _GEN_1457;
  assign rf_matrix_b_4_tile_v_3_MPORT_14_addr = 8'h61;
  assign rf_matrix_b_4_tile_v_3_MPORT_14_data = rf[rf_matrix_b_4_tile_v_3_MPORT_14_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_4_tile_v_2_MPORT_14_en = handshaked & _GEN_1457;
  assign rf_matrix_b_4_tile_v_2_MPORT_14_addr = 8'h65;
  assign rf_matrix_b_4_tile_v_2_MPORT_14_data = rf[rf_matrix_b_4_tile_v_2_MPORT_14_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_4_tile_v_1_MPORT_14_en = handshaked & _GEN_1457;
  assign rf_matrix_b_4_tile_v_1_MPORT_14_addr = 8'h69;
  assign rf_matrix_b_4_tile_v_1_MPORT_14_data = rf[rf_matrix_b_4_tile_v_1_MPORT_14_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_4_tile_v_0_MPORT_14_en = handshaked & _GEN_1457;
  assign rf_matrix_b_4_tile_v_0_MPORT_14_addr = 8'h6d;
  assign rf_matrix_b_4_tile_v_0_MPORT_14_data = rf[rf_matrix_b_4_tile_v_0_MPORT_14_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_4_tile_v_3_MPORT_14_en = handshaked & _GEN_1457;
  assign rf_matrix_c_4_tile_v_3_MPORT_14_addr = 8'hb0;
  assign rf_matrix_c_4_tile_v_3_MPORT_14_data = rf[rf_matrix_c_4_tile_v_3_MPORT_14_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_4_tile_v_2_MPORT_14_en = handshaked & _GEN_1457;
  assign rf_matrix_c_4_tile_v_2_MPORT_14_addr = 8'hb1;
  assign rf_matrix_c_4_tile_v_2_MPORT_14_data = rf[rf_matrix_c_4_tile_v_2_MPORT_14_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_4_tile_v_1_MPORT_14_en = handshaked & _GEN_1457;
  assign rf_matrix_c_4_tile_v_1_MPORT_14_addr = 8'hb8;
  assign rf_matrix_c_4_tile_v_1_MPORT_14_data = rf[rf_matrix_c_4_tile_v_1_MPORT_14_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_4_tile_v_0_MPORT_14_en = handshaked & _GEN_1457;
  assign rf_matrix_c_4_tile_v_0_MPORT_14_addr = 8'hb9;
  assign rf_matrix_c_4_tile_v_0_MPORT_14_data = rf[rf_matrix_c_4_tile_v_0_MPORT_14_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_3_MPORT_37_en = handshaked & _GEN_1469;
  assign rf_a_tile_v_3_MPORT_37_addr = 8'h12;
  assign rf_a_tile_v_3_MPORT_37_data = rf[rf_a_tile_v_3_MPORT_37_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_2_MPORT_37_en = handshaked & _GEN_1469;
  assign rf_a_tile_v_2_MPORT_37_addr = 8'h16;
  assign rf_a_tile_v_2_MPORT_37_data = rf[rf_a_tile_v_2_MPORT_37_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_1_MPORT_111_en = handshaked & _GEN_1469;
  assign rf_a_tile_v_1_MPORT_111_addr = 8'h1a;
  assign rf_a_tile_v_1_MPORT_111_data = rf[rf_a_tile_v_1_MPORT_111_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_0_MPORT_111_en = handshaked & _GEN_1469;
  assign rf_a_tile_v_0_MPORT_111_addr = 8'h1e;
  assign rf_a_tile_v_0_MPORT_111_data = rf[rf_a_tile_v_0_MPORT_111_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_4_tile_v_3_MPORT_15_en = handshaked & _GEN_1469;
  assign rf_matrix_b_4_tile_v_3_MPORT_15_addr = 8'h61;
  assign rf_matrix_b_4_tile_v_3_MPORT_15_data = rf[rf_matrix_b_4_tile_v_3_MPORT_15_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_4_tile_v_2_MPORT_15_en = handshaked & _GEN_1469;
  assign rf_matrix_b_4_tile_v_2_MPORT_15_addr = 8'h65;
  assign rf_matrix_b_4_tile_v_2_MPORT_15_data = rf[rf_matrix_b_4_tile_v_2_MPORT_15_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_4_tile_v_1_MPORT_15_en = handshaked & _GEN_1469;
  assign rf_matrix_b_4_tile_v_1_MPORT_15_addr = 8'h69;
  assign rf_matrix_b_4_tile_v_1_MPORT_15_data = rf[rf_matrix_b_4_tile_v_1_MPORT_15_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_4_tile_v_0_MPORT_15_en = handshaked & _GEN_1469;
  assign rf_matrix_b_4_tile_v_0_MPORT_15_addr = 8'h6d;
  assign rf_matrix_b_4_tile_v_0_MPORT_15_data = rf[rf_matrix_b_4_tile_v_0_MPORT_15_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_4_tile_v_3_MPORT_15_en = handshaked & _GEN_1469;
  assign rf_matrix_c_4_tile_v_3_MPORT_15_addr = 8'h91;
  assign rf_matrix_c_4_tile_v_3_MPORT_15_data = rf[rf_matrix_c_4_tile_v_3_MPORT_15_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_4_tile_v_2_MPORT_15_en = handshaked & _GEN_1469;
  assign rf_matrix_c_4_tile_v_2_MPORT_15_addr = 8'h95;
  assign rf_matrix_c_4_tile_v_2_MPORT_15_data = rf[rf_matrix_c_4_tile_v_2_MPORT_15_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_4_tile_v_1_MPORT_15_en = handshaked & _GEN_1469;
  assign rf_matrix_c_4_tile_v_1_MPORT_15_addr = 8'h99;
  assign rf_matrix_c_4_tile_v_1_MPORT_15_data = rf[rf_matrix_c_4_tile_v_1_MPORT_15_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_4_tile_v_0_MPORT_15_en = handshaked & _GEN_1469;
  assign rf_matrix_c_4_tile_v_0_MPORT_15_addr = 8'h9d;
  assign rf_matrix_c_4_tile_v_0_MPORT_15_data = rf[rf_matrix_c_4_tile_v_0_MPORT_15_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_1_MPORT_112_en = handshaked & _GEN_1483;
  assign rf_a_tile_v_1_MPORT_112_addr = 8'h12;
  assign rf_a_tile_v_1_MPORT_112_data = rf[rf_a_tile_v_1_MPORT_112_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_0_MPORT_112_en = handshaked & _GEN_1483;
  assign rf_a_tile_v_0_MPORT_112_addr = 8'h16;
  assign rf_a_tile_v_0_MPORT_112_data = rf[rf_a_tile_v_0_MPORT_112_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_4_tile_v_3_MPORT_16_en = handshaked & _GEN_1483;
  assign rf_matrix_b_4_tile_v_3_MPORT_16_addr = 8'h61;
  assign rf_matrix_b_4_tile_v_3_MPORT_16_data = rf[rf_matrix_b_4_tile_v_3_MPORT_16_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_4_tile_v_2_MPORT_16_en = handshaked & _GEN_1483;
  assign rf_matrix_b_4_tile_v_2_MPORT_16_addr = 8'h65;
  assign rf_matrix_b_4_tile_v_2_MPORT_16_data = rf[rf_matrix_b_4_tile_v_2_MPORT_16_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_4_tile_v_1_MPORT_16_en = handshaked & _GEN_1483;
  assign rf_matrix_b_4_tile_v_1_MPORT_16_addr = 8'h69;
  assign rf_matrix_b_4_tile_v_1_MPORT_16_data = rf[rf_matrix_b_4_tile_v_1_MPORT_16_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_4_tile_v_0_MPORT_16_en = handshaked & _GEN_1483;
  assign rf_matrix_b_4_tile_v_0_MPORT_16_addr = 8'h6d;
  assign rf_matrix_b_4_tile_v_0_MPORT_16_data = rf[rf_matrix_b_4_tile_v_0_MPORT_16_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_4_tile_v_3_MPORT_16_en = handshaked & _GEN_1483;
  assign rf_matrix_c_4_tile_v_3_MPORT_16_addr = 8'ha2;
  assign rf_matrix_c_4_tile_v_3_MPORT_16_data = rf[rf_matrix_c_4_tile_v_3_MPORT_16_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_4_tile_v_2_MPORT_16_en = handshaked & _GEN_1483;
  assign rf_matrix_c_4_tile_v_2_MPORT_16_addr = 8'ha3;
  assign rf_matrix_c_4_tile_v_2_MPORT_16_data = rf[rf_matrix_c_4_tile_v_2_MPORT_16_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_4_tile_v_1_MPORT_16_en = handshaked & _GEN_1483;
  assign rf_matrix_c_4_tile_v_1_MPORT_16_addr = 8'haa;
  assign rf_matrix_c_4_tile_v_1_MPORT_16_data = rf[rf_matrix_c_4_tile_v_1_MPORT_16_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_4_tile_v_0_MPORT_16_en = handshaked & _GEN_1483;
  assign rf_matrix_c_4_tile_v_0_MPORT_16_addr = 8'hab;
  assign rf_matrix_c_4_tile_v_0_MPORT_16_data = rf[rf_matrix_c_4_tile_v_0_MPORT_16_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_1_MPORT_113_en = handshaked & _GEN_1495;
  assign rf_a_tile_v_1_MPORT_113_addr = 8'h1a;
  assign rf_a_tile_v_1_MPORT_113_data = rf[rf_a_tile_v_1_MPORT_113_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_0_MPORT_113_en = handshaked & _GEN_1495;
  assign rf_a_tile_v_0_MPORT_113_addr = 8'h1e;
  assign rf_a_tile_v_0_MPORT_113_data = rf[rf_a_tile_v_0_MPORT_113_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_4_tile_v_3_MPORT_17_en = handshaked & _GEN_1495;
  assign rf_matrix_b_4_tile_v_3_MPORT_17_addr = 8'h61;
  assign rf_matrix_b_4_tile_v_3_MPORT_17_data = rf[rf_matrix_b_4_tile_v_3_MPORT_17_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_4_tile_v_2_MPORT_17_en = handshaked & _GEN_1495;
  assign rf_matrix_b_4_tile_v_2_MPORT_17_addr = 8'h65;
  assign rf_matrix_b_4_tile_v_2_MPORT_17_data = rf[rf_matrix_b_4_tile_v_2_MPORT_17_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_4_tile_v_1_MPORT_17_en = handshaked & _GEN_1495;
  assign rf_matrix_b_4_tile_v_1_MPORT_17_addr = 8'h69;
  assign rf_matrix_b_4_tile_v_1_MPORT_17_data = rf[rf_matrix_b_4_tile_v_1_MPORT_17_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_4_tile_v_0_MPORT_17_en = handshaked & _GEN_1495;
  assign rf_matrix_b_4_tile_v_0_MPORT_17_addr = 8'h6d;
  assign rf_matrix_b_4_tile_v_0_MPORT_17_data = rf[rf_matrix_b_4_tile_v_0_MPORT_17_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_4_tile_v_3_MPORT_17_en = handshaked & _GEN_1495;
  assign rf_matrix_c_4_tile_v_3_MPORT_17_addr = 8'hb2;
  assign rf_matrix_c_4_tile_v_3_MPORT_17_data = rf[rf_matrix_c_4_tile_v_3_MPORT_17_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_4_tile_v_2_MPORT_17_en = handshaked & _GEN_1495;
  assign rf_matrix_c_4_tile_v_2_MPORT_17_addr = 8'hb3;
  assign rf_matrix_c_4_tile_v_2_MPORT_17_data = rf[rf_matrix_c_4_tile_v_2_MPORT_17_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_4_tile_v_1_MPORT_17_en = handshaked & _GEN_1495;
  assign rf_matrix_c_4_tile_v_1_MPORT_17_addr = 8'hba;
  assign rf_matrix_c_4_tile_v_1_MPORT_17_data = rf[rf_matrix_c_4_tile_v_1_MPORT_17_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_4_tile_v_0_MPORT_17_en = handshaked & _GEN_1495;
  assign rf_matrix_c_4_tile_v_0_MPORT_17_addr = 8'hbb;
  assign rf_matrix_c_4_tile_v_0_MPORT_17_data = rf[rf_matrix_c_4_tile_v_0_MPORT_17_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_1_MPORT_114_en = handshaked & _GEN_1507;
  assign rf_a_tile_v_1_MPORT_114_addr = 8'h13;
  assign rf_a_tile_v_1_MPORT_114_data = rf[rf_a_tile_v_1_MPORT_114_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_0_MPORT_114_en = handshaked & _GEN_1507;
  assign rf_a_tile_v_0_MPORT_114_addr = 8'h17;
  assign rf_a_tile_v_0_MPORT_114_data = rf[rf_a_tile_v_0_MPORT_114_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_4_tile_v_3_MPORT_18_en = handshaked & _GEN_1507;
  assign rf_matrix_b_4_tile_v_3_MPORT_18_addr = 8'h71;
  assign rf_matrix_b_4_tile_v_3_MPORT_18_data = rf[rf_matrix_b_4_tile_v_3_MPORT_18_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_4_tile_v_2_MPORT_18_en = handshaked & _GEN_1507;
  assign rf_matrix_b_4_tile_v_2_MPORT_18_addr = 8'h75;
  assign rf_matrix_b_4_tile_v_2_MPORT_18_data = rf[rf_matrix_b_4_tile_v_2_MPORT_18_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_4_tile_v_1_MPORT_18_en = handshaked & _GEN_1507;
  assign rf_matrix_b_4_tile_v_1_MPORT_18_addr = 8'h79;
  assign rf_matrix_b_4_tile_v_1_MPORT_18_data = rf[rf_matrix_b_4_tile_v_1_MPORT_18_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_4_tile_v_0_MPORT_18_en = handshaked & _GEN_1507;
  assign rf_matrix_b_4_tile_v_0_MPORT_18_addr = 8'h7d;
  assign rf_matrix_b_4_tile_v_0_MPORT_18_data = rf[rf_matrix_b_4_tile_v_0_MPORT_18_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_4_tile_v_3_MPORT_18_en = handshaked & _GEN_1507;
  assign rf_matrix_c_4_tile_v_3_MPORT_18_addr = 8'ha0;
  assign rf_matrix_c_4_tile_v_3_MPORT_18_data = rf[rf_matrix_c_4_tile_v_3_MPORT_18_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_4_tile_v_2_MPORT_18_en = handshaked & _GEN_1507;
  assign rf_matrix_c_4_tile_v_2_MPORT_18_addr = 8'ha1;
  assign rf_matrix_c_4_tile_v_2_MPORT_18_data = rf[rf_matrix_c_4_tile_v_2_MPORT_18_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_4_tile_v_1_MPORT_18_en = handshaked & _GEN_1507;
  assign rf_matrix_c_4_tile_v_1_MPORT_18_addr = 8'ha8;
  assign rf_matrix_c_4_tile_v_1_MPORT_18_data = rf[rf_matrix_c_4_tile_v_1_MPORT_18_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_4_tile_v_0_MPORT_18_en = handshaked & _GEN_1507;
  assign rf_matrix_c_4_tile_v_0_MPORT_18_addr = 8'ha9;
  assign rf_matrix_c_4_tile_v_0_MPORT_18_data = rf[rf_matrix_c_4_tile_v_0_MPORT_18_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_3_MPORT_38_en = handshaked & _GEN_1519;
  assign rf_a_tile_v_3_MPORT_38_addr = 8'h13;
  assign rf_a_tile_v_3_MPORT_38_data = rf[rf_a_tile_v_3_MPORT_38_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_2_MPORT_38_en = handshaked & _GEN_1519;
  assign rf_a_tile_v_2_MPORT_38_addr = 8'h17;
  assign rf_a_tile_v_2_MPORT_38_data = rf[rf_a_tile_v_2_MPORT_38_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_1_MPORT_115_en = handshaked & _GEN_1519;
  assign rf_a_tile_v_1_MPORT_115_addr = 8'h1b;
  assign rf_a_tile_v_1_MPORT_115_data = rf[rf_a_tile_v_1_MPORT_115_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_0_MPORT_115_en = handshaked & _GEN_1519;
  assign rf_a_tile_v_0_MPORT_115_addr = 8'h1f;
  assign rf_a_tile_v_0_MPORT_115_data = rf[rf_a_tile_v_0_MPORT_115_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_4_tile_v_3_MPORT_19_en = handshaked & _GEN_1519;
  assign rf_matrix_b_4_tile_v_3_MPORT_19_addr = 8'h71;
  assign rf_matrix_b_4_tile_v_3_MPORT_19_data = rf[rf_matrix_b_4_tile_v_3_MPORT_19_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_4_tile_v_2_MPORT_19_en = handshaked & _GEN_1519;
  assign rf_matrix_b_4_tile_v_2_MPORT_19_addr = 8'h75;
  assign rf_matrix_b_4_tile_v_2_MPORT_19_data = rf[rf_matrix_b_4_tile_v_2_MPORT_19_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_4_tile_v_1_MPORT_19_en = handshaked & _GEN_1519;
  assign rf_matrix_b_4_tile_v_1_MPORT_19_addr = 8'h79;
  assign rf_matrix_b_4_tile_v_1_MPORT_19_data = rf[rf_matrix_b_4_tile_v_1_MPORT_19_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_4_tile_v_0_MPORT_19_en = handshaked & _GEN_1519;
  assign rf_matrix_b_4_tile_v_0_MPORT_19_addr = 8'h7d;
  assign rf_matrix_b_4_tile_v_0_MPORT_19_data = rf[rf_matrix_b_4_tile_v_0_MPORT_19_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_4_tile_v_3_MPORT_19_en = handshaked & _GEN_1519;
  assign rf_matrix_c_4_tile_v_3_MPORT_19_addr = 8'h90;
  assign rf_matrix_c_4_tile_v_3_MPORT_19_data = rf[rf_matrix_c_4_tile_v_3_MPORT_19_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_4_tile_v_2_MPORT_19_en = handshaked & _GEN_1519;
  assign rf_matrix_c_4_tile_v_2_MPORT_19_addr = 8'h94;
  assign rf_matrix_c_4_tile_v_2_MPORT_19_data = rf[rf_matrix_c_4_tile_v_2_MPORT_19_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_4_tile_v_1_MPORT_19_en = handshaked & _GEN_1519;
  assign rf_matrix_c_4_tile_v_1_MPORT_19_addr = 8'h98;
  assign rf_matrix_c_4_tile_v_1_MPORT_19_data = rf[rf_matrix_c_4_tile_v_1_MPORT_19_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_4_tile_v_0_MPORT_19_en = handshaked & _GEN_1519;
  assign rf_matrix_c_4_tile_v_0_MPORT_19_addr = 8'h9c;
  assign rf_matrix_c_4_tile_v_0_MPORT_19_data = rf[rf_matrix_c_4_tile_v_0_MPORT_19_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_1_MPORT_116_en = handshaked & _GEN_1533;
  assign rf_a_tile_v_1_MPORT_116_addr = 8'h1b;
  assign rf_a_tile_v_1_MPORT_116_data = rf[rf_a_tile_v_1_MPORT_116_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_0_MPORT_116_en = handshaked & _GEN_1533;
  assign rf_a_tile_v_0_MPORT_116_addr = 8'h1f;
  assign rf_a_tile_v_0_MPORT_116_data = rf[rf_a_tile_v_0_MPORT_116_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_4_tile_v_3_MPORT_20_en = handshaked & _GEN_1533;
  assign rf_matrix_b_4_tile_v_3_MPORT_20_addr = 8'h71;
  assign rf_matrix_b_4_tile_v_3_MPORT_20_data = rf[rf_matrix_b_4_tile_v_3_MPORT_20_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_4_tile_v_2_MPORT_20_en = handshaked & _GEN_1533;
  assign rf_matrix_b_4_tile_v_2_MPORT_20_addr = 8'h75;
  assign rf_matrix_b_4_tile_v_2_MPORT_20_data = rf[rf_matrix_b_4_tile_v_2_MPORT_20_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_4_tile_v_1_MPORT_20_en = handshaked & _GEN_1533;
  assign rf_matrix_b_4_tile_v_1_MPORT_20_addr = 8'h79;
  assign rf_matrix_b_4_tile_v_1_MPORT_20_data = rf[rf_matrix_b_4_tile_v_1_MPORT_20_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_4_tile_v_0_MPORT_20_en = handshaked & _GEN_1533;
  assign rf_matrix_b_4_tile_v_0_MPORT_20_addr = 8'h7d;
  assign rf_matrix_b_4_tile_v_0_MPORT_20_data = rf[rf_matrix_b_4_tile_v_0_MPORT_20_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_4_tile_v_3_MPORT_20_en = handshaked & _GEN_1533;
  assign rf_matrix_c_4_tile_v_3_MPORT_20_addr = 8'hb0;
  assign rf_matrix_c_4_tile_v_3_MPORT_20_data = rf[rf_matrix_c_4_tile_v_3_MPORT_20_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_4_tile_v_2_MPORT_20_en = handshaked & _GEN_1533;
  assign rf_matrix_c_4_tile_v_2_MPORT_20_addr = 8'hb1;
  assign rf_matrix_c_4_tile_v_2_MPORT_20_data = rf[rf_matrix_c_4_tile_v_2_MPORT_20_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_4_tile_v_1_MPORT_20_en = handshaked & _GEN_1533;
  assign rf_matrix_c_4_tile_v_1_MPORT_20_addr = 8'hb8;
  assign rf_matrix_c_4_tile_v_1_MPORT_20_data = rf[rf_matrix_c_4_tile_v_1_MPORT_20_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_4_tile_v_0_MPORT_20_en = handshaked & _GEN_1533;
  assign rf_matrix_c_4_tile_v_0_MPORT_20_addr = 8'hb9;
  assign rf_matrix_c_4_tile_v_0_MPORT_20_data = rf[rf_matrix_c_4_tile_v_0_MPORT_20_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_3_MPORT_39_en = handshaked & _GEN_1545;
  assign rf_a_tile_v_3_MPORT_39_addr = 8'h13;
  assign rf_a_tile_v_3_MPORT_39_data = rf[rf_a_tile_v_3_MPORT_39_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_2_MPORT_39_en = handshaked & _GEN_1545;
  assign rf_a_tile_v_2_MPORT_39_addr = 8'h17;
  assign rf_a_tile_v_2_MPORT_39_data = rf[rf_a_tile_v_2_MPORT_39_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_1_MPORT_117_en = handshaked & _GEN_1545;
  assign rf_a_tile_v_1_MPORT_117_addr = 8'h1b;
  assign rf_a_tile_v_1_MPORT_117_data = rf[rf_a_tile_v_1_MPORT_117_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_0_MPORT_117_en = handshaked & _GEN_1545;
  assign rf_a_tile_v_0_MPORT_117_addr = 8'h1f;
  assign rf_a_tile_v_0_MPORT_117_data = rf[rf_a_tile_v_0_MPORT_117_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_4_tile_v_3_MPORT_21_en = handshaked & _GEN_1545;
  assign rf_matrix_b_4_tile_v_3_MPORT_21_addr = 8'h71;
  assign rf_matrix_b_4_tile_v_3_MPORT_21_data = rf[rf_matrix_b_4_tile_v_3_MPORT_21_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_4_tile_v_2_MPORT_21_en = handshaked & _GEN_1545;
  assign rf_matrix_b_4_tile_v_2_MPORT_21_addr = 8'h75;
  assign rf_matrix_b_4_tile_v_2_MPORT_21_data = rf[rf_matrix_b_4_tile_v_2_MPORT_21_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_4_tile_v_1_MPORT_21_en = handshaked & _GEN_1545;
  assign rf_matrix_b_4_tile_v_1_MPORT_21_addr = 8'h79;
  assign rf_matrix_b_4_tile_v_1_MPORT_21_data = rf[rf_matrix_b_4_tile_v_1_MPORT_21_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_4_tile_v_0_MPORT_21_en = handshaked & _GEN_1545;
  assign rf_matrix_b_4_tile_v_0_MPORT_21_addr = 8'h7d;
  assign rf_matrix_b_4_tile_v_0_MPORT_21_data = rf[rf_matrix_b_4_tile_v_0_MPORT_21_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_4_tile_v_3_MPORT_21_en = handshaked & _GEN_1545;
  assign rf_matrix_c_4_tile_v_3_MPORT_21_addr = 8'h91;
  assign rf_matrix_c_4_tile_v_3_MPORT_21_data = rf[rf_matrix_c_4_tile_v_3_MPORT_21_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_4_tile_v_2_MPORT_21_en = handshaked & _GEN_1545;
  assign rf_matrix_c_4_tile_v_2_MPORT_21_addr = 8'h95;
  assign rf_matrix_c_4_tile_v_2_MPORT_21_data = rf[rf_matrix_c_4_tile_v_2_MPORT_21_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_4_tile_v_1_MPORT_21_en = handshaked & _GEN_1545;
  assign rf_matrix_c_4_tile_v_1_MPORT_21_addr = 8'h99;
  assign rf_matrix_c_4_tile_v_1_MPORT_21_data = rf[rf_matrix_c_4_tile_v_1_MPORT_21_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_4_tile_v_0_MPORT_21_en = handshaked & _GEN_1545;
  assign rf_matrix_c_4_tile_v_0_MPORT_21_addr = 8'h9d;
  assign rf_matrix_c_4_tile_v_0_MPORT_21_data = rf[rf_matrix_c_4_tile_v_0_MPORT_21_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_1_MPORT_118_en = handshaked & _GEN_1559;
  assign rf_a_tile_v_1_MPORT_118_addr = 8'h13;
  assign rf_a_tile_v_1_MPORT_118_data = rf[rf_a_tile_v_1_MPORT_118_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_0_MPORT_118_en = handshaked & _GEN_1559;
  assign rf_a_tile_v_0_MPORT_118_addr = 8'h17;
  assign rf_a_tile_v_0_MPORT_118_data = rf[rf_a_tile_v_0_MPORT_118_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_4_tile_v_3_MPORT_22_en = handshaked & _GEN_1559;
  assign rf_matrix_b_4_tile_v_3_MPORT_22_addr = 8'h71;
  assign rf_matrix_b_4_tile_v_3_MPORT_22_data = rf[rf_matrix_b_4_tile_v_3_MPORT_22_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_4_tile_v_2_MPORT_22_en = handshaked & _GEN_1559;
  assign rf_matrix_b_4_tile_v_2_MPORT_22_addr = 8'h75;
  assign rf_matrix_b_4_tile_v_2_MPORT_22_data = rf[rf_matrix_b_4_tile_v_2_MPORT_22_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_4_tile_v_1_MPORT_22_en = handshaked & _GEN_1559;
  assign rf_matrix_b_4_tile_v_1_MPORT_22_addr = 8'h79;
  assign rf_matrix_b_4_tile_v_1_MPORT_22_data = rf[rf_matrix_b_4_tile_v_1_MPORT_22_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_4_tile_v_0_MPORT_22_en = handshaked & _GEN_1559;
  assign rf_matrix_b_4_tile_v_0_MPORT_22_addr = 8'h7d;
  assign rf_matrix_b_4_tile_v_0_MPORT_22_data = rf[rf_matrix_b_4_tile_v_0_MPORT_22_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_4_tile_v_3_MPORT_22_en = handshaked & _GEN_1559;
  assign rf_matrix_c_4_tile_v_3_MPORT_22_addr = 8'ha2;
  assign rf_matrix_c_4_tile_v_3_MPORT_22_data = rf[rf_matrix_c_4_tile_v_3_MPORT_22_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_4_tile_v_2_MPORT_22_en = handshaked & _GEN_1559;
  assign rf_matrix_c_4_tile_v_2_MPORT_22_addr = 8'ha3;
  assign rf_matrix_c_4_tile_v_2_MPORT_22_data = rf[rf_matrix_c_4_tile_v_2_MPORT_22_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_4_tile_v_1_MPORT_22_en = handshaked & _GEN_1559;
  assign rf_matrix_c_4_tile_v_1_MPORT_22_addr = 8'haa;
  assign rf_matrix_c_4_tile_v_1_MPORT_22_data = rf[rf_matrix_c_4_tile_v_1_MPORT_22_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_4_tile_v_0_MPORT_22_en = handshaked & _GEN_1559;
  assign rf_matrix_c_4_tile_v_0_MPORT_22_addr = 8'hab;
  assign rf_matrix_c_4_tile_v_0_MPORT_22_data = rf[rf_matrix_c_4_tile_v_0_MPORT_22_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_1_MPORT_119_en = handshaked & _GEN_1571;
  assign rf_a_tile_v_1_MPORT_119_addr = 8'h1b;
  assign rf_a_tile_v_1_MPORT_119_data = rf[rf_a_tile_v_1_MPORT_119_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_0_MPORT_119_en = handshaked & _GEN_1571;
  assign rf_a_tile_v_0_MPORT_119_addr = 8'h1f;
  assign rf_a_tile_v_0_MPORT_119_data = rf[rf_a_tile_v_0_MPORT_119_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_4_tile_v_3_MPORT_23_en = handshaked & _GEN_1571;
  assign rf_matrix_b_4_tile_v_3_MPORT_23_addr = 8'h71;
  assign rf_matrix_b_4_tile_v_3_MPORT_23_data = rf[rf_matrix_b_4_tile_v_3_MPORT_23_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_4_tile_v_2_MPORT_23_en = handshaked & _GEN_1571;
  assign rf_matrix_b_4_tile_v_2_MPORT_23_addr = 8'h75;
  assign rf_matrix_b_4_tile_v_2_MPORT_23_data = rf[rf_matrix_b_4_tile_v_2_MPORT_23_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_4_tile_v_1_MPORT_23_en = handshaked & _GEN_1571;
  assign rf_matrix_b_4_tile_v_1_MPORT_23_addr = 8'h79;
  assign rf_matrix_b_4_tile_v_1_MPORT_23_data = rf[rf_matrix_b_4_tile_v_1_MPORT_23_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_4_tile_v_0_MPORT_23_en = handshaked & _GEN_1571;
  assign rf_matrix_b_4_tile_v_0_MPORT_23_addr = 8'h7d;
  assign rf_matrix_b_4_tile_v_0_MPORT_23_data = rf[rf_matrix_b_4_tile_v_0_MPORT_23_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_4_tile_v_3_MPORT_23_en = handshaked & _GEN_1571;
  assign rf_matrix_c_4_tile_v_3_MPORT_23_addr = 8'hb2;
  assign rf_matrix_c_4_tile_v_3_MPORT_23_data = rf[rf_matrix_c_4_tile_v_3_MPORT_23_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_4_tile_v_2_MPORT_23_en = handshaked & _GEN_1571;
  assign rf_matrix_c_4_tile_v_2_MPORT_23_addr = 8'hb3;
  assign rf_matrix_c_4_tile_v_2_MPORT_23_data = rf[rf_matrix_c_4_tile_v_2_MPORT_23_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_4_tile_v_1_MPORT_23_en = handshaked & _GEN_1571;
  assign rf_matrix_c_4_tile_v_1_MPORT_23_addr = 8'hba;
  assign rf_matrix_c_4_tile_v_1_MPORT_23_data = rf[rf_matrix_c_4_tile_v_1_MPORT_23_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_4_tile_v_0_MPORT_23_en = handshaked & _GEN_1571;
  assign rf_matrix_c_4_tile_v_0_MPORT_23_addr = 8'hbb;
  assign rf_matrix_c_4_tile_v_0_MPORT_23_data = rf[rf_matrix_c_4_tile_v_0_MPORT_23_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_1_MPORT_120_en = handshaked & _GEN_1276;
  assign rf_a_tile_v_1_MPORT_120_addr = 8'h30;
  assign rf_a_tile_v_1_MPORT_120_data = rf[rf_a_tile_v_1_MPORT_120_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_0_MPORT_120_en = handshaked & _GEN_1276;
  assign rf_a_tile_v_0_MPORT_120_addr = 8'h34;
  assign rf_a_tile_v_0_MPORT_120_data = rf[rf_a_tile_v_0_MPORT_120_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_5_tile_v_3_MPORT_en = handshaked & _GEN_1276;
  assign rf_matrix_b_5_tile_v_3_MPORT_addr = 8'h41;
  assign rf_matrix_b_5_tile_v_3_MPORT_data = rf[rf_matrix_b_5_tile_v_3_MPORT_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_5_tile_v_2_MPORT_en = handshaked & _GEN_1276;
  assign rf_matrix_b_5_tile_v_2_MPORT_addr = 8'h45;
  assign rf_matrix_b_5_tile_v_2_MPORT_data = rf[rf_matrix_b_5_tile_v_2_MPORT_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_5_tile_v_1_MPORT_en = handshaked & _GEN_1276;
  assign rf_matrix_b_5_tile_v_1_MPORT_addr = 8'h49;
  assign rf_matrix_b_5_tile_v_1_MPORT_data = rf[rf_matrix_b_5_tile_v_1_MPORT_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_5_tile_v_0_MPORT_en = handshaked & _GEN_1276;
  assign rf_matrix_b_5_tile_v_0_MPORT_addr = 8'h4d;
  assign rf_matrix_b_5_tile_v_0_MPORT_data = rf[rf_matrix_b_5_tile_v_0_MPORT_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_5_tile_v_3_MPORT_en = handshaked & _GEN_1276;
  assign rf_matrix_c_5_tile_v_3_MPORT_addr = 8'he0;
  assign rf_matrix_c_5_tile_v_3_MPORT_data = rf[rf_matrix_c_5_tile_v_3_MPORT_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_5_tile_v_2_MPORT_en = handshaked & _GEN_1276;
  assign rf_matrix_c_5_tile_v_2_MPORT_addr = 8'he1;
  assign rf_matrix_c_5_tile_v_2_MPORT_data = rf[rf_matrix_c_5_tile_v_2_MPORT_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_5_tile_v_1_MPORT_en = handshaked & _GEN_1276;
  assign rf_matrix_c_5_tile_v_1_MPORT_addr = 8'he8;
  assign rf_matrix_c_5_tile_v_1_MPORT_data = rf[rf_matrix_c_5_tile_v_1_MPORT_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_5_tile_v_0_MPORT_en = handshaked & _GEN_1276;
  assign rf_matrix_c_5_tile_v_0_MPORT_addr = 8'he9;
  assign rf_matrix_c_5_tile_v_0_MPORT_data = rf[rf_matrix_c_5_tile_v_0_MPORT_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_3_MPORT_40_en = handshaked & _GEN_1291;
  assign rf_a_tile_v_3_MPORT_40_addr = 8'h30;
  assign rf_a_tile_v_3_MPORT_40_data = rf[rf_a_tile_v_3_MPORT_40_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_2_MPORT_40_en = handshaked & _GEN_1291;
  assign rf_a_tile_v_2_MPORT_40_addr = 8'h34;
  assign rf_a_tile_v_2_MPORT_40_data = rf[rf_a_tile_v_2_MPORT_40_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_1_MPORT_121_en = handshaked & _GEN_1291;
  assign rf_a_tile_v_1_MPORT_121_addr = 8'h38;
  assign rf_a_tile_v_1_MPORT_121_data = rf[rf_a_tile_v_1_MPORT_121_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_0_MPORT_121_en = handshaked & _GEN_1291;
  assign rf_a_tile_v_0_MPORT_121_addr = 8'h3c;
  assign rf_a_tile_v_0_MPORT_121_data = rf[rf_a_tile_v_0_MPORT_121_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_5_tile_v_3_MPORT_1_en = handshaked & _GEN_1291;
  assign rf_matrix_b_5_tile_v_3_MPORT_1_addr = 8'h41;
  assign rf_matrix_b_5_tile_v_3_MPORT_1_data = rf[rf_matrix_b_5_tile_v_3_MPORT_1_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_5_tile_v_2_MPORT_1_en = handshaked & _GEN_1291;
  assign rf_matrix_b_5_tile_v_2_MPORT_1_addr = 8'h45;
  assign rf_matrix_b_5_tile_v_2_MPORT_1_data = rf[rf_matrix_b_5_tile_v_2_MPORT_1_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_5_tile_v_1_MPORT_1_en = handshaked & _GEN_1291;
  assign rf_matrix_b_5_tile_v_1_MPORT_1_addr = 8'h49;
  assign rf_matrix_b_5_tile_v_1_MPORT_1_data = rf[rf_matrix_b_5_tile_v_1_MPORT_1_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_5_tile_v_0_MPORT_1_en = handshaked & _GEN_1291;
  assign rf_matrix_b_5_tile_v_0_MPORT_1_addr = 8'h4d;
  assign rf_matrix_b_5_tile_v_0_MPORT_1_data = rf[rf_matrix_b_5_tile_v_0_MPORT_1_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_5_tile_v_3_MPORT_1_en = handshaked & _GEN_1291;
  assign rf_matrix_c_5_tile_v_3_MPORT_1_addr = 8'hb0;
  assign rf_matrix_c_5_tile_v_3_MPORT_1_data = rf[rf_matrix_c_5_tile_v_3_MPORT_1_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_5_tile_v_2_MPORT_1_en = handshaked & _GEN_1291;
  assign rf_matrix_c_5_tile_v_2_MPORT_1_addr = 8'hb4;
  assign rf_matrix_c_5_tile_v_2_MPORT_1_data = rf[rf_matrix_c_5_tile_v_2_MPORT_1_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_5_tile_v_1_MPORT_1_en = handshaked & _GEN_1291;
  assign rf_matrix_c_5_tile_v_1_MPORT_1_addr = 8'hb8;
  assign rf_matrix_c_5_tile_v_1_MPORT_1_data = rf[rf_matrix_c_5_tile_v_1_MPORT_1_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_5_tile_v_0_MPORT_1_en = handshaked & _GEN_1291;
  assign rf_matrix_c_5_tile_v_0_MPORT_1_addr = 8'hbc;
  assign rf_matrix_c_5_tile_v_0_MPORT_1_data = rf[rf_matrix_c_5_tile_v_0_MPORT_1_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_1_MPORT_122_en = handshaked & _GEN_1305;
  assign rf_a_tile_v_1_MPORT_122_addr = 8'h38;
  assign rf_a_tile_v_1_MPORT_122_data = rf[rf_a_tile_v_1_MPORT_122_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_0_MPORT_122_en = handshaked & _GEN_1305;
  assign rf_a_tile_v_0_MPORT_122_addr = 8'h3c;
  assign rf_a_tile_v_0_MPORT_122_data = rf[rf_a_tile_v_0_MPORT_122_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_5_tile_v_3_MPORT_2_en = handshaked & _GEN_1305;
  assign rf_matrix_b_5_tile_v_3_MPORT_2_addr = 8'h41;
  assign rf_matrix_b_5_tile_v_3_MPORT_2_data = rf[rf_matrix_b_5_tile_v_3_MPORT_2_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_5_tile_v_2_MPORT_2_en = handshaked & _GEN_1305;
  assign rf_matrix_b_5_tile_v_2_MPORT_2_addr = 8'h45;
  assign rf_matrix_b_5_tile_v_2_MPORT_2_data = rf[rf_matrix_b_5_tile_v_2_MPORT_2_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_5_tile_v_1_MPORT_2_en = handshaked & _GEN_1305;
  assign rf_matrix_b_5_tile_v_1_MPORT_2_addr = 8'h49;
  assign rf_matrix_b_5_tile_v_1_MPORT_2_data = rf[rf_matrix_b_5_tile_v_1_MPORT_2_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_5_tile_v_0_MPORT_2_en = handshaked & _GEN_1305;
  assign rf_matrix_b_5_tile_v_0_MPORT_2_addr = 8'h4d;
  assign rf_matrix_b_5_tile_v_0_MPORT_2_data = rf[rf_matrix_b_5_tile_v_0_MPORT_2_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_5_tile_v_3_MPORT_2_en = handshaked & _GEN_1305;
  assign rf_matrix_c_5_tile_v_3_MPORT_2_addr = 8'hf0;
  assign rf_matrix_c_5_tile_v_3_MPORT_2_data = rf[rf_matrix_c_5_tile_v_3_MPORT_2_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_5_tile_v_2_MPORT_2_en = handshaked & _GEN_1305;
  assign rf_matrix_c_5_tile_v_2_MPORT_2_addr = 8'hf1;
  assign rf_matrix_c_5_tile_v_2_MPORT_2_data = rf[rf_matrix_c_5_tile_v_2_MPORT_2_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_5_tile_v_1_MPORT_2_en = handshaked & _GEN_1305;
  assign rf_matrix_c_5_tile_v_1_MPORT_2_addr = 8'hf8;
  assign rf_matrix_c_5_tile_v_1_MPORT_2_data = rf[rf_matrix_c_5_tile_v_1_MPORT_2_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_5_tile_v_0_MPORT_2_en = handshaked & _GEN_1305;
  assign rf_matrix_c_5_tile_v_0_MPORT_2_addr = 8'hf9;
  assign rf_matrix_c_5_tile_v_0_MPORT_2_data = rf[rf_matrix_c_5_tile_v_0_MPORT_2_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_3_MPORT_41_en = handshaked & _GEN_1317;
  assign rf_a_tile_v_3_MPORT_41_addr = 8'h30;
  assign rf_a_tile_v_3_MPORT_41_data = rf[rf_a_tile_v_3_MPORT_41_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_2_MPORT_41_en = handshaked & _GEN_1317;
  assign rf_a_tile_v_2_MPORT_41_addr = 8'h34;
  assign rf_a_tile_v_2_MPORT_41_data = rf[rf_a_tile_v_2_MPORT_41_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_1_MPORT_123_en = handshaked & _GEN_1317;
  assign rf_a_tile_v_1_MPORT_123_addr = 8'h38;
  assign rf_a_tile_v_1_MPORT_123_data = rf[rf_a_tile_v_1_MPORT_123_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_0_MPORT_123_en = handshaked & _GEN_1317;
  assign rf_a_tile_v_0_MPORT_123_addr = 8'h3c;
  assign rf_a_tile_v_0_MPORT_123_data = rf[rf_a_tile_v_0_MPORT_123_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_5_tile_v_3_MPORT_3_en = handshaked & _GEN_1317;
  assign rf_matrix_b_5_tile_v_3_MPORT_3_addr = 8'h41;
  assign rf_matrix_b_5_tile_v_3_MPORT_3_data = rf[rf_matrix_b_5_tile_v_3_MPORT_3_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_5_tile_v_2_MPORT_3_en = handshaked & _GEN_1317;
  assign rf_matrix_b_5_tile_v_2_MPORT_3_addr = 8'h45;
  assign rf_matrix_b_5_tile_v_2_MPORT_3_data = rf[rf_matrix_b_5_tile_v_2_MPORT_3_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_5_tile_v_1_MPORT_3_en = handshaked & _GEN_1317;
  assign rf_matrix_b_5_tile_v_1_MPORT_3_addr = 8'h49;
  assign rf_matrix_b_5_tile_v_1_MPORT_3_data = rf[rf_matrix_b_5_tile_v_1_MPORT_3_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_5_tile_v_0_MPORT_3_en = handshaked & _GEN_1317;
  assign rf_matrix_b_5_tile_v_0_MPORT_3_addr = 8'h4d;
  assign rf_matrix_b_5_tile_v_0_MPORT_3_data = rf[rf_matrix_b_5_tile_v_0_MPORT_3_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_5_tile_v_3_MPORT_3_en = handshaked & _GEN_1317;
  assign rf_matrix_c_5_tile_v_3_MPORT_3_addr = 8'hb1;
  assign rf_matrix_c_5_tile_v_3_MPORT_3_data = rf[rf_matrix_c_5_tile_v_3_MPORT_3_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_5_tile_v_2_MPORT_3_en = handshaked & _GEN_1317;
  assign rf_matrix_c_5_tile_v_2_MPORT_3_addr = 8'hb5;
  assign rf_matrix_c_5_tile_v_2_MPORT_3_data = rf[rf_matrix_c_5_tile_v_2_MPORT_3_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_5_tile_v_1_MPORT_3_en = handshaked & _GEN_1317;
  assign rf_matrix_c_5_tile_v_1_MPORT_3_addr = 8'hb9;
  assign rf_matrix_c_5_tile_v_1_MPORT_3_data = rf[rf_matrix_c_5_tile_v_1_MPORT_3_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_5_tile_v_0_MPORT_3_en = handshaked & _GEN_1317;
  assign rf_matrix_c_5_tile_v_0_MPORT_3_addr = 8'hbd;
  assign rf_matrix_c_5_tile_v_0_MPORT_3_data = rf[rf_matrix_c_5_tile_v_0_MPORT_3_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_1_MPORT_124_en = handshaked & _GEN_1331;
  assign rf_a_tile_v_1_MPORT_124_addr = 8'h30;
  assign rf_a_tile_v_1_MPORT_124_data = rf[rf_a_tile_v_1_MPORT_124_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_0_MPORT_124_en = handshaked & _GEN_1331;
  assign rf_a_tile_v_0_MPORT_124_addr = 8'h34;
  assign rf_a_tile_v_0_MPORT_124_data = rf[rf_a_tile_v_0_MPORT_124_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_5_tile_v_3_MPORT_4_en = handshaked & _GEN_1331;
  assign rf_matrix_b_5_tile_v_3_MPORT_4_addr = 8'h41;
  assign rf_matrix_b_5_tile_v_3_MPORT_4_data = rf[rf_matrix_b_5_tile_v_3_MPORT_4_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_5_tile_v_2_MPORT_4_en = handshaked & _GEN_1331;
  assign rf_matrix_b_5_tile_v_2_MPORT_4_addr = 8'h45;
  assign rf_matrix_b_5_tile_v_2_MPORT_4_data = rf[rf_matrix_b_5_tile_v_2_MPORT_4_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_5_tile_v_1_MPORT_4_en = handshaked & _GEN_1331;
  assign rf_matrix_b_5_tile_v_1_MPORT_4_addr = 8'h49;
  assign rf_matrix_b_5_tile_v_1_MPORT_4_data = rf[rf_matrix_b_5_tile_v_1_MPORT_4_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_5_tile_v_0_MPORT_4_en = handshaked & _GEN_1331;
  assign rf_matrix_b_5_tile_v_0_MPORT_4_addr = 8'h4d;
  assign rf_matrix_b_5_tile_v_0_MPORT_4_data = rf[rf_matrix_b_5_tile_v_0_MPORT_4_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_5_tile_v_3_MPORT_4_en = handshaked & _GEN_1331;
  assign rf_matrix_c_5_tile_v_3_MPORT_4_addr = 8'he2;
  assign rf_matrix_c_5_tile_v_3_MPORT_4_data = rf[rf_matrix_c_5_tile_v_3_MPORT_4_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_5_tile_v_2_MPORT_4_en = handshaked & _GEN_1331;
  assign rf_matrix_c_5_tile_v_2_MPORT_4_addr = 8'he3;
  assign rf_matrix_c_5_tile_v_2_MPORT_4_data = rf[rf_matrix_c_5_tile_v_2_MPORT_4_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_5_tile_v_1_MPORT_4_en = handshaked & _GEN_1331;
  assign rf_matrix_c_5_tile_v_1_MPORT_4_addr = 8'hea;
  assign rf_matrix_c_5_tile_v_1_MPORT_4_data = rf[rf_matrix_c_5_tile_v_1_MPORT_4_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_5_tile_v_0_MPORT_4_en = handshaked & _GEN_1331;
  assign rf_matrix_c_5_tile_v_0_MPORT_4_addr = 8'heb;
  assign rf_matrix_c_5_tile_v_0_MPORT_4_data = rf[rf_matrix_c_5_tile_v_0_MPORT_4_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_1_MPORT_125_en = handshaked & _GEN_1343;
  assign rf_a_tile_v_1_MPORT_125_addr = 8'h38;
  assign rf_a_tile_v_1_MPORT_125_data = rf[rf_a_tile_v_1_MPORT_125_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_0_MPORT_125_en = handshaked & _GEN_1343;
  assign rf_a_tile_v_0_MPORT_125_addr = 8'h3c;
  assign rf_a_tile_v_0_MPORT_125_data = rf[rf_a_tile_v_0_MPORT_125_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_5_tile_v_3_MPORT_5_en = handshaked & _GEN_1343;
  assign rf_matrix_b_5_tile_v_3_MPORT_5_addr = 8'h41;
  assign rf_matrix_b_5_tile_v_3_MPORT_5_data = rf[rf_matrix_b_5_tile_v_3_MPORT_5_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_5_tile_v_2_MPORT_5_en = handshaked & _GEN_1343;
  assign rf_matrix_b_5_tile_v_2_MPORT_5_addr = 8'h45;
  assign rf_matrix_b_5_tile_v_2_MPORT_5_data = rf[rf_matrix_b_5_tile_v_2_MPORT_5_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_5_tile_v_1_MPORT_5_en = handshaked & _GEN_1343;
  assign rf_matrix_b_5_tile_v_1_MPORT_5_addr = 8'h49;
  assign rf_matrix_b_5_tile_v_1_MPORT_5_data = rf[rf_matrix_b_5_tile_v_1_MPORT_5_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_5_tile_v_0_MPORT_5_en = handshaked & _GEN_1343;
  assign rf_matrix_b_5_tile_v_0_MPORT_5_addr = 8'h4d;
  assign rf_matrix_b_5_tile_v_0_MPORT_5_data = rf[rf_matrix_b_5_tile_v_0_MPORT_5_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_5_tile_v_3_MPORT_5_en = handshaked & _GEN_1343;
  assign rf_matrix_c_5_tile_v_3_MPORT_5_addr = 8'hf2;
  assign rf_matrix_c_5_tile_v_3_MPORT_5_data = rf[rf_matrix_c_5_tile_v_3_MPORT_5_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_5_tile_v_2_MPORT_5_en = handshaked & _GEN_1343;
  assign rf_matrix_c_5_tile_v_2_MPORT_5_addr = 8'hf3;
  assign rf_matrix_c_5_tile_v_2_MPORT_5_data = rf[rf_matrix_c_5_tile_v_2_MPORT_5_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_5_tile_v_1_MPORT_5_en = handshaked & _GEN_1343;
  assign rf_matrix_c_5_tile_v_1_MPORT_5_addr = 8'hfa;
  assign rf_matrix_c_5_tile_v_1_MPORT_5_data = rf[rf_matrix_c_5_tile_v_1_MPORT_5_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_5_tile_v_0_MPORT_5_en = handshaked & _GEN_1343;
  assign rf_matrix_c_5_tile_v_0_MPORT_5_addr = 8'hfb;
  assign rf_matrix_c_5_tile_v_0_MPORT_5_data = rf[rf_matrix_c_5_tile_v_0_MPORT_5_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_1_MPORT_126_en = handshaked & _GEN_1355;
  assign rf_a_tile_v_1_MPORT_126_addr = 8'h31;
  assign rf_a_tile_v_1_MPORT_126_data = rf[rf_a_tile_v_1_MPORT_126_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_0_MPORT_126_en = handshaked & _GEN_1355;
  assign rf_a_tile_v_0_MPORT_126_addr = 8'h35;
  assign rf_a_tile_v_0_MPORT_126_data = rf[rf_a_tile_v_0_MPORT_126_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_5_tile_v_3_MPORT_6_en = handshaked & _GEN_1355;
  assign rf_matrix_b_5_tile_v_3_MPORT_6_addr = 8'h51;
  assign rf_matrix_b_5_tile_v_3_MPORT_6_data = rf[rf_matrix_b_5_tile_v_3_MPORT_6_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_5_tile_v_2_MPORT_6_en = handshaked & _GEN_1355;
  assign rf_matrix_b_5_tile_v_2_MPORT_6_addr = 8'h55;
  assign rf_matrix_b_5_tile_v_2_MPORT_6_data = rf[rf_matrix_b_5_tile_v_2_MPORT_6_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_5_tile_v_1_MPORT_6_en = handshaked & _GEN_1355;
  assign rf_matrix_b_5_tile_v_1_MPORT_6_addr = 8'h59;
  assign rf_matrix_b_5_tile_v_1_MPORT_6_data = rf[rf_matrix_b_5_tile_v_1_MPORT_6_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_5_tile_v_0_MPORT_6_en = handshaked & _GEN_1355;
  assign rf_matrix_b_5_tile_v_0_MPORT_6_addr = 8'h5d;
  assign rf_matrix_b_5_tile_v_0_MPORT_6_data = rf[rf_matrix_b_5_tile_v_0_MPORT_6_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_5_tile_v_3_MPORT_6_en = handshaked & _GEN_1355;
  assign rf_matrix_c_5_tile_v_3_MPORT_6_addr = 8'he0;
  assign rf_matrix_c_5_tile_v_3_MPORT_6_data = rf[rf_matrix_c_5_tile_v_3_MPORT_6_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_5_tile_v_2_MPORT_6_en = handshaked & _GEN_1355;
  assign rf_matrix_c_5_tile_v_2_MPORT_6_addr = 8'he1;
  assign rf_matrix_c_5_tile_v_2_MPORT_6_data = rf[rf_matrix_c_5_tile_v_2_MPORT_6_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_5_tile_v_1_MPORT_6_en = handshaked & _GEN_1355;
  assign rf_matrix_c_5_tile_v_1_MPORT_6_addr = 8'he8;
  assign rf_matrix_c_5_tile_v_1_MPORT_6_data = rf[rf_matrix_c_5_tile_v_1_MPORT_6_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_5_tile_v_0_MPORT_6_en = handshaked & _GEN_1355;
  assign rf_matrix_c_5_tile_v_0_MPORT_6_addr = 8'he9;
  assign rf_matrix_c_5_tile_v_0_MPORT_6_data = rf[rf_matrix_c_5_tile_v_0_MPORT_6_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_3_MPORT_42_en = handshaked & _GEN_1367;
  assign rf_a_tile_v_3_MPORT_42_addr = 8'h31;
  assign rf_a_tile_v_3_MPORT_42_data = rf[rf_a_tile_v_3_MPORT_42_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_2_MPORT_42_en = handshaked & _GEN_1367;
  assign rf_a_tile_v_2_MPORT_42_addr = 8'h35;
  assign rf_a_tile_v_2_MPORT_42_data = rf[rf_a_tile_v_2_MPORT_42_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_1_MPORT_127_en = handshaked & _GEN_1367;
  assign rf_a_tile_v_1_MPORT_127_addr = 8'h39;
  assign rf_a_tile_v_1_MPORT_127_data = rf[rf_a_tile_v_1_MPORT_127_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_0_MPORT_127_en = handshaked & _GEN_1367;
  assign rf_a_tile_v_0_MPORT_127_addr = 8'h3d;
  assign rf_a_tile_v_0_MPORT_127_data = rf[rf_a_tile_v_0_MPORT_127_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_5_tile_v_3_MPORT_7_en = handshaked & _GEN_1367;
  assign rf_matrix_b_5_tile_v_3_MPORT_7_addr = 8'h51;
  assign rf_matrix_b_5_tile_v_3_MPORT_7_data = rf[rf_matrix_b_5_tile_v_3_MPORT_7_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_5_tile_v_2_MPORT_7_en = handshaked & _GEN_1367;
  assign rf_matrix_b_5_tile_v_2_MPORT_7_addr = 8'h55;
  assign rf_matrix_b_5_tile_v_2_MPORT_7_data = rf[rf_matrix_b_5_tile_v_2_MPORT_7_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_5_tile_v_1_MPORT_7_en = handshaked & _GEN_1367;
  assign rf_matrix_b_5_tile_v_1_MPORT_7_addr = 8'h59;
  assign rf_matrix_b_5_tile_v_1_MPORT_7_data = rf[rf_matrix_b_5_tile_v_1_MPORT_7_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_5_tile_v_0_MPORT_7_en = handshaked & _GEN_1367;
  assign rf_matrix_b_5_tile_v_0_MPORT_7_addr = 8'h5d;
  assign rf_matrix_b_5_tile_v_0_MPORT_7_data = rf[rf_matrix_b_5_tile_v_0_MPORT_7_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_5_tile_v_3_MPORT_7_en = handshaked & _GEN_1367;
  assign rf_matrix_c_5_tile_v_3_MPORT_7_addr = 8'hb0;
  assign rf_matrix_c_5_tile_v_3_MPORT_7_data = rf[rf_matrix_c_5_tile_v_3_MPORT_7_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_5_tile_v_2_MPORT_7_en = handshaked & _GEN_1367;
  assign rf_matrix_c_5_tile_v_2_MPORT_7_addr = 8'hb4;
  assign rf_matrix_c_5_tile_v_2_MPORT_7_data = rf[rf_matrix_c_5_tile_v_2_MPORT_7_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_5_tile_v_1_MPORT_7_en = handshaked & _GEN_1367;
  assign rf_matrix_c_5_tile_v_1_MPORT_7_addr = 8'hb8;
  assign rf_matrix_c_5_tile_v_1_MPORT_7_data = rf[rf_matrix_c_5_tile_v_1_MPORT_7_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_5_tile_v_0_MPORT_7_en = handshaked & _GEN_1367;
  assign rf_matrix_c_5_tile_v_0_MPORT_7_addr = 8'hbc;
  assign rf_matrix_c_5_tile_v_0_MPORT_7_data = rf[rf_matrix_c_5_tile_v_0_MPORT_7_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_1_MPORT_128_en = handshaked & _GEN_1381;
  assign rf_a_tile_v_1_MPORT_128_addr = 8'h39;
  assign rf_a_tile_v_1_MPORT_128_data = rf[rf_a_tile_v_1_MPORT_128_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_0_MPORT_128_en = handshaked & _GEN_1381;
  assign rf_a_tile_v_0_MPORT_128_addr = 8'h3d;
  assign rf_a_tile_v_0_MPORT_128_data = rf[rf_a_tile_v_0_MPORT_128_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_5_tile_v_3_MPORT_8_en = handshaked & _GEN_1381;
  assign rf_matrix_b_5_tile_v_3_MPORT_8_addr = 8'h51;
  assign rf_matrix_b_5_tile_v_3_MPORT_8_data = rf[rf_matrix_b_5_tile_v_3_MPORT_8_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_5_tile_v_2_MPORT_8_en = handshaked & _GEN_1381;
  assign rf_matrix_b_5_tile_v_2_MPORT_8_addr = 8'h55;
  assign rf_matrix_b_5_tile_v_2_MPORT_8_data = rf[rf_matrix_b_5_tile_v_2_MPORT_8_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_5_tile_v_1_MPORT_8_en = handshaked & _GEN_1381;
  assign rf_matrix_b_5_tile_v_1_MPORT_8_addr = 8'h59;
  assign rf_matrix_b_5_tile_v_1_MPORT_8_data = rf[rf_matrix_b_5_tile_v_1_MPORT_8_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_5_tile_v_0_MPORT_8_en = handshaked & _GEN_1381;
  assign rf_matrix_b_5_tile_v_0_MPORT_8_addr = 8'h5d;
  assign rf_matrix_b_5_tile_v_0_MPORT_8_data = rf[rf_matrix_b_5_tile_v_0_MPORT_8_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_5_tile_v_3_MPORT_8_en = handshaked & _GEN_1381;
  assign rf_matrix_c_5_tile_v_3_MPORT_8_addr = 8'hf0;
  assign rf_matrix_c_5_tile_v_3_MPORT_8_data = rf[rf_matrix_c_5_tile_v_3_MPORT_8_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_5_tile_v_2_MPORT_8_en = handshaked & _GEN_1381;
  assign rf_matrix_c_5_tile_v_2_MPORT_8_addr = 8'hf1;
  assign rf_matrix_c_5_tile_v_2_MPORT_8_data = rf[rf_matrix_c_5_tile_v_2_MPORT_8_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_5_tile_v_1_MPORT_8_en = handshaked & _GEN_1381;
  assign rf_matrix_c_5_tile_v_1_MPORT_8_addr = 8'hf8;
  assign rf_matrix_c_5_tile_v_1_MPORT_8_data = rf[rf_matrix_c_5_tile_v_1_MPORT_8_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_5_tile_v_0_MPORT_8_en = handshaked & _GEN_1381;
  assign rf_matrix_c_5_tile_v_0_MPORT_8_addr = 8'hf9;
  assign rf_matrix_c_5_tile_v_0_MPORT_8_data = rf[rf_matrix_c_5_tile_v_0_MPORT_8_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_3_MPORT_43_en = handshaked & _GEN_1393;
  assign rf_a_tile_v_3_MPORT_43_addr = 8'h31;
  assign rf_a_tile_v_3_MPORT_43_data = rf[rf_a_tile_v_3_MPORT_43_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_2_MPORT_43_en = handshaked & _GEN_1393;
  assign rf_a_tile_v_2_MPORT_43_addr = 8'h35;
  assign rf_a_tile_v_2_MPORT_43_data = rf[rf_a_tile_v_2_MPORT_43_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_1_MPORT_129_en = handshaked & _GEN_1393;
  assign rf_a_tile_v_1_MPORT_129_addr = 8'h39;
  assign rf_a_tile_v_1_MPORT_129_data = rf[rf_a_tile_v_1_MPORT_129_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_0_MPORT_129_en = handshaked & _GEN_1393;
  assign rf_a_tile_v_0_MPORT_129_addr = 8'h3d;
  assign rf_a_tile_v_0_MPORT_129_data = rf[rf_a_tile_v_0_MPORT_129_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_5_tile_v_3_MPORT_9_en = handshaked & _GEN_1393;
  assign rf_matrix_b_5_tile_v_3_MPORT_9_addr = 8'h51;
  assign rf_matrix_b_5_tile_v_3_MPORT_9_data = rf[rf_matrix_b_5_tile_v_3_MPORT_9_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_5_tile_v_2_MPORT_9_en = handshaked & _GEN_1393;
  assign rf_matrix_b_5_tile_v_2_MPORT_9_addr = 8'h55;
  assign rf_matrix_b_5_tile_v_2_MPORT_9_data = rf[rf_matrix_b_5_tile_v_2_MPORT_9_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_5_tile_v_1_MPORT_9_en = handshaked & _GEN_1393;
  assign rf_matrix_b_5_tile_v_1_MPORT_9_addr = 8'h59;
  assign rf_matrix_b_5_tile_v_1_MPORT_9_data = rf[rf_matrix_b_5_tile_v_1_MPORT_9_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_5_tile_v_0_MPORT_9_en = handshaked & _GEN_1393;
  assign rf_matrix_b_5_tile_v_0_MPORT_9_addr = 8'h5d;
  assign rf_matrix_b_5_tile_v_0_MPORT_9_data = rf[rf_matrix_b_5_tile_v_0_MPORT_9_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_5_tile_v_3_MPORT_9_en = handshaked & _GEN_1393;
  assign rf_matrix_c_5_tile_v_3_MPORT_9_addr = 8'hb1;
  assign rf_matrix_c_5_tile_v_3_MPORT_9_data = rf[rf_matrix_c_5_tile_v_3_MPORT_9_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_5_tile_v_2_MPORT_9_en = handshaked & _GEN_1393;
  assign rf_matrix_c_5_tile_v_2_MPORT_9_addr = 8'hb5;
  assign rf_matrix_c_5_tile_v_2_MPORT_9_data = rf[rf_matrix_c_5_tile_v_2_MPORT_9_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_5_tile_v_1_MPORT_9_en = handshaked & _GEN_1393;
  assign rf_matrix_c_5_tile_v_1_MPORT_9_addr = 8'hb9;
  assign rf_matrix_c_5_tile_v_1_MPORT_9_data = rf[rf_matrix_c_5_tile_v_1_MPORT_9_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_5_tile_v_0_MPORT_9_en = handshaked & _GEN_1393;
  assign rf_matrix_c_5_tile_v_0_MPORT_9_addr = 8'hbd;
  assign rf_matrix_c_5_tile_v_0_MPORT_9_data = rf[rf_matrix_c_5_tile_v_0_MPORT_9_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_1_MPORT_130_en = handshaked & _GEN_1407;
  assign rf_a_tile_v_1_MPORT_130_addr = 8'h31;
  assign rf_a_tile_v_1_MPORT_130_data = rf[rf_a_tile_v_1_MPORT_130_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_0_MPORT_130_en = handshaked & _GEN_1407;
  assign rf_a_tile_v_0_MPORT_130_addr = 8'h35;
  assign rf_a_tile_v_0_MPORT_130_data = rf[rf_a_tile_v_0_MPORT_130_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_5_tile_v_3_MPORT_10_en = handshaked & _GEN_1407;
  assign rf_matrix_b_5_tile_v_3_MPORT_10_addr = 8'h51;
  assign rf_matrix_b_5_tile_v_3_MPORT_10_data = rf[rf_matrix_b_5_tile_v_3_MPORT_10_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_5_tile_v_2_MPORT_10_en = handshaked & _GEN_1407;
  assign rf_matrix_b_5_tile_v_2_MPORT_10_addr = 8'h55;
  assign rf_matrix_b_5_tile_v_2_MPORT_10_data = rf[rf_matrix_b_5_tile_v_2_MPORT_10_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_5_tile_v_1_MPORT_10_en = handshaked & _GEN_1407;
  assign rf_matrix_b_5_tile_v_1_MPORT_10_addr = 8'h59;
  assign rf_matrix_b_5_tile_v_1_MPORT_10_data = rf[rf_matrix_b_5_tile_v_1_MPORT_10_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_5_tile_v_0_MPORT_10_en = handshaked & _GEN_1407;
  assign rf_matrix_b_5_tile_v_0_MPORT_10_addr = 8'h5d;
  assign rf_matrix_b_5_tile_v_0_MPORT_10_data = rf[rf_matrix_b_5_tile_v_0_MPORT_10_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_5_tile_v_3_MPORT_10_en = handshaked & _GEN_1407;
  assign rf_matrix_c_5_tile_v_3_MPORT_10_addr = 8'he2;
  assign rf_matrix_c_5_tile_v_3_MPORT_10_data = rf[rf_matrix_c_5_tile_v_3_MPORT_10_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_5_tile_v_2_MPORT_10_en = handshaked & _GEN_1407;
  assign rf_matrix_c_5_tile_v_2_MPORT_10_addr = 8'he3;
  assign rf_matrix_c_5_tile_v_2_MPORT_10_data = rf[rf_matrix_c_5_tile_v_2_MPORT_10_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_5_tile_v_1_MPORT_10_en = handshaked & _GEN_1407;
  assign rf_matrix_c_5_tile_v_1_MPORT_10_addr = 8'hea;
  assign rf_matrix_c_5_tile_v_1_MPORT_10_data = rf[rf_matrix_c_5_tile_v_1_MPORT_10_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_5_tile_v_0_MPORT_10_en = handshaked & _GEN_1407;
  assign rf_matrix_c_5_tile_v_0_MPORT_10_addr = 8'heb;
  assign rf_matrix_c_5_tile_v_0_MPORT_10_data = rf[rf_matrix_c_5_tile_v_0_MPORT_10_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_1_MPORT_131_en = handshaked & _GEN_1419;
  assign rf_a_tile_v_1_MPORT_131_addr = 8'h39;
  assign rf_a_tile_v_1_MPORT_131_data = rf[rf_a_tile_v_1_MPORT_131_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_0_MPORT_131_en = handshaked & _GEN_1419;
  assign rf_a_tile_v_0_MPORT_131_addr = 8'h3d;
  assign rf_a_tile_v_0_MPORT_131_data = rf[rf_a_tile_v_0_MPORT_131_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_5_tile_v_3_MPORT_11_en = handshaked & _GEN_1419;
  assign rf_matrix_b_5_tile_v_3_MPORT_11_addr = 8'h51;
  assign rf_matrix_b_5_tile_v_3_MPORT_11_data = rf[rf_matrix_b_5_tile_v_3_MPORT_11_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_5_tile_v_2_MPORT_11_en = handshaked & _GEN_1419;
  assign rf_matrix_b_5_tile_v_2_MPORT_11_addr = 8'h55;
  assign rf_matrix_b_5_tile_v_2_MPORT_11_data = rf[rf_matrix_b_5_tile_v_2_MPORT_11_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_5_tile_v_1_MPORT_11_en = handshaked & _GEN_1419;
  assign rf_matrix_b_5_tile_v_1_MPORT_11_addr = 8'h59;
  assign rf_matrix_b_5_tile_v_1_MPORT_11_data = rf[rf_matrix_b_5_tile_v_1_MPORT_11_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_5_tile_v_0_MPORT_11_en = handshaked & _GEN_1419;
  assign rf_matrix_b_5_tile_v_0_MPORT_11_addr = 8'h5d;
  assign rf_matrix_b_5_tile_v_0_MPORT_11_data = rf[rf_matrix_b_5_tile_v_0_MPORT_11_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_5_tile_v_3_MPORT_11_en = handshaked & _GEN_1419;
  assign rf_matrix_c_5_tile_v_3_MPORT_11_addr = 8'hf2;
  assign rf_matrix_c_5_tile_v_3_MPORT_11_data = rf[rf_matrix_c_5_tile_v_3_MPORT_11_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_5_tile_v_2_MPORT_11_en = handshaked & _GEN_1419;
  assign rf_matrix_c_5_tile_v_2_MPORT_11_addr = 8'hf3;
  assign rf_matrix_c_5_tile_v_2_MPORT_11_data = rf[rf_matrix_c_5_tile_v_2_MPORT_11_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_5_tile_v_1_MPORT_11_en = handshaked & _GEN_1419;
  assign rf_matrix_c_5_tile_v_1_MPORT_11_addr = 8'hfa;
  assign rf_matrix_c_5_tile_v_1_MPORT_11_data = rf[rf_matrix_c_5_tile_v_1_MPORT_11_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_5_tile_v_0_MPORT_11_en = handshaked & _GEN_1419;
  assign rf_matrix_c_5_tile_v_0_MPORT_11_addr = 8'hfb;
  assign rf_matrix_c_5_tile_v_0_MPORT_11_data = rf[rf_matrix_c_5_tile_v_0_MPORT_11_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_1_MPORT_132_en = handshaked & _GEN_1431;
  assign rf_a_tile_v_1_MPORT_132_addr = 8'h32;
  assign rf_a_tile_v_1_MPORT_132_data = rf[rf_a_tile_v_1_MPORT_132_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_0_MPORT_132_en = handshaked & _GEN_1431;
  assign rf_a_tile_v_0_MPORT_132_addr = 8'h36;
  assign rf_a_tile_v_0_MPORT_132_data = rf[rf_a_tile_v_0_MPORT_132_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_5_tile_v_3_MPORT_12_en = handshaked & _GEN_1431;
  assign rf_matrix_b_5_tile_v_3_MPORT_12_addr = 8'h61;
  assign rf_matrix_b_5_tile_v_3_MPORT_12_data = rf[rf_matrix_b_5_tile_v_3_MPORT_12_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_5_tile_v_2_MPORT_12_en = handshaked & _GEN_1431;
  assign rf_matrix_b_5_tile_v_2_MPORT_12_addr = 8'h65;
  assign rf_matrix_b_5_tile_v_2_MPORT_12_data = rf[rf_matrix_b_5_tile_v_2_MPORT_12_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_5_tile_v_1_MPORT_12_en = handshaked & _GEN_1431;
  assign rf_matrix_b_5_tile_v_1_MPORT_12_addr = 8'h69;
  assign rf_matrix_b_5_tile_v_1_MPORT_12_data = rf[rf_matrix_b_5_tile_v_1_MPORT_12_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_5_tile_v_0_MPORT_12_en = handshaked & _GEN_1431;
  assign rf_matrix_b_5_tile_v_0_MPORT_12_addr = 8'h6d;
  assign rf_matrix_b_5_tile_v_0_MPORT_12_data = rf[rf_matrix_b_5_tile_v_0_MPORT_12_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_5_tile_v_3_MPORT_12_en = handshaked & _GEN_1431;
  assign rf_matrix_c_5_tile_v_3_MPORT_12_addr = 8'he0;
  assign rf_matrix_c_5_tile_v_3_MPORT_12_data = rf[rf_matrix_c_5_tile_v_3_MPORT_12_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_5_tile_v_2_MPORT_12_en = handshaked & _GEN_1431;
  assign rf_matrix_c_5_tile_v_2_MPORT_12_addr = 8'he1;
  assign rf_matrix_c_5_tile_v_2_MPORT_12_data = rf[rf_matrix_c_5_tile_v_2_MPORT_12_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_5_tile_v_1_MPORT_12_en = handshaked & _GEN_1431;
  assign rf_matrix_c_5_tile_v_1_MPORT_12_addr = 8'he8;
  assign rf_matrix_c_5_tile_v_1_MPORT_12_data = rf[rf_matrix_c_5_tile_v_1_MPORT_12_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_5_tile_v_0_MPORT_12_en = handshaked & _GEN_1431;
  assign rf_matrix_c_5_tile_v_0_MPORT_12_addr = 8'he9;
  assign rf_matrix_c_5_tile_v_0_MPORT_12_data = rf[rf_matrix_c_5_tile_v_0_MPORT_12_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_3_MPORT_44_en = handshaked & _GEN_1443;
  assign rf_a_tile_v_3_MPORT_44_addr = 8'h32;
  assign rf_a_tile_v_3_MPORT_44_data = rf[rf_a_tile_v_3_MPORT_44_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_2_MPORT_44_en = handshaked & _GEN_1443;
  assign rf_a_tile_v_2_MPORT_44_addr = 8'h36;
  assign rf_a_tile_v_2_MPORT_44_data = rf[rf_a_tile_v_2_MPORT_44_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_1_MPORT_133_en = handshaked & _GEN_1443;
  assign rf_a_tile_v_1_MPORT_133_addr = 8'h3a;
  assign rf_a_tile_v_1_MPORT_133_data = rf[rf_a_tile_v_1_MPORT_133_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_0_MPORT_133_en = handshaked & _GEN_1443;
  assign rf_a_tile_v_0_MPORT_133_addr = 8'h3e;
  assign rf_a_tile_v_0_MPORT_133_data = rf[rf_a_tile_v_0_MPORT_133_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_5_tile_v_3_MPORT_13_en = handshaked & _GEN_1443;
  assign rf_matrix_b_5_tile_v_3_MPORT_13_addr = 8'h61;
  assign rf_matrix_b_5_tile_v_3_MPORT_13_data = rf[rf_matrix_b_5_tile_v_3_MPORT_13_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_5_tile_v_2_MPORT_13_en = handshaked & _GEN_1443;
  assign rf_matrix_b_5_tile_v_2_MPORT_13_addr = 8'h65;
  assign rf_matrix_b_5_tile_v_2_MPORT_13_data = rf[rf_matrix_b_5_tile_v_2_MPORT_13_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_5_tile_v_1_MPORT_13_en = handshaked & _GEN_1443;
  assign rf_matrix_b_5_tile_v_1_MPORT_13_addr = 8'h69;
  assign rf_matrix_b_5_tile_v_1_MPORT_13_data = rf[rf_matrix_b_5_tile_v_1_MPORT_13_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_5_tile_v_0_MPORT_13_en = handshaked & _GEN_1443;
  assign rf_matrix_b_5_tile_v_0_MPORT_13_addr = 8'h6d;
  assign rf_matrix_b_5_tile_v_0_MPORT_13_data = rf[rf_matrix_b_5_tile_v_0_MPORT_13_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_5_tile_v_3_MPORT_13_en = handshaked & _GEN_1443;
  assign rf_matrix_c_5_tile_v_3_MPORT_13_addr = 8'hb0;
  assign rf_matrix_c_5_tile_v_3_MPORT_13_data = rf[rf_matrix_c_5_tile_v_3_MPORT_13_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_5_tile_v_2_MPORT_13_en = handshaked & _GEN_1443;
  assign rf_matrix_c_5_tile_v_2_MPORT_13_addr = 8'hb4;
  assign rf_matrix_c_5_tile_v_2_MPORT_13_data = rf[rf_matrix_c_5_tile_v_2_MPORT_13_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_5_tile_v_1_MPORT_13_en = handshaked & _GEN_1443;
  assign rf_matrix_c_5_tile_v_1_MPORT_13_addr = 8'hb8;
  assign rf_matrix_c_5_tile_v_1_MPORT_13_data = rf[rf_matrix_c_5_tile_v_1_MPORT_13_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_5_tile_v_0_MPORT_13_en = handshaked & _GEN_1443;
  assign rf_matrix_c_5_tile_v_0_MPORT_13_addr = 8'hbc;
  assign rf_matrix_c_5_tile_v_0_MPORT_13_data = rf[rf_matrix_c_5_tile_v_0_MPORT_13_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_1_MPORT_134_en = handshaked & _GEN_1457;
  assign rf_a_tile_v_1_MPORT_134_addr = 8'h3a;
  assign rf_a_tile_v_1_MPORT_134_data = rf[rf_a_tile_v_1_MPORT_134_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_0_MPORT_134_en = handshaked & _GEN_1457;
  assign rf_a_tile_v_0_MPORT_134_addr = 8'h3e;
  assign rf_a_tile_v_0_MPORT_134_data = rf[rf_a_tile_v_0_MPORT_134_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_5_tile_v_3_MPORT_14_en = handshaked & _GEN_1457;
  assign rf_matrix_b_5_tile_v_3_MPORT_14_addr = 8'h61;
  assign rf_matrix_b_5_tile_v_3_MPORT_14_data = rf[rf_matrix_b_5_tile_v_3_MPORT_14_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_5_tile_v_2_MPORT_14_en = handshaked & _GEN_1457;
  assign rf_matrix_b_5_tile_v_2_MPORT_14_addr = 8'h65;
  assign rf_matrix_b_5_tile_v_2_MPORT_14_data = rf[rf_matrix_b_5_tile_v_2_MPORT_14_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_5_tile_v_1_MPORT_14_en = handshaked & _GEN_1457;
  assign rf_matrix_b_5_tile_v_1_MPORT_14_addr = 8'h69;
  assign rf_matrix_b_5_tile_v_1_MPORT_14_data = rf[rf_matrix_b_5_tile_v_1_MPORT_14_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_5_tile_v_0_MPORT_14_en = handshaked & _GEN_1457;
  assign rf_matrix_b_5_tile_v_0_MPORT_14_addr = 8'h6d;
  assign rf_matrix_b_5_tile_v_0_MPORT_14_data = rf[rf_matrix_b_5_tile_v_0_MPORT_14_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_5_tile_v_3_MPORT_14_en = handshaked & _GEN_1457;
  assign rf_matrix_c_5_tile_v_3_MPORT_14_addr = 8'hf0;
  assign rf_matrix_c_5_tile_v_3_MPORT_14_data = rf[rf_matrix_c_5_tile_v_3_MPORT_14_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_5_tile_v_2_MPORT_14_en = handshaked & _GEN_1457;
  assign rf_matrix_c_5_tile_v_2_MPORT_14_addr = 8'hf1;
  assign rf_matrix_c_5_tile_v_2_MPORT_14_data = rf[rf_matrix_c_5_tile_v_2_MPORT_14_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_5_tile_v_1_MPORT_14_en = handshaked & _GEN_1457;
  assign rf_matrix_c_5_tile_v_1_MPORT_14_addr = 8'hf8;
  assign rf_matrix_c_5_tile_v_1_MPORT_14_data = rf[rf_matrix_c_5_tile_v_1_MPORT_14_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_5_tile_v_0_MPORT_14_en = handshaked & _GEN_1457;
  assign rf_matrix_c_5_tile_v_0_MPORT_14_addr = 8'hf9;
  assign rf_matrix_c_5_tile_v_0_MPORT_14_data = rf[rf_matrix_c_5_tile_v_0_MPORT_14_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_3_MPORT_45_en = handshaked & _GEN_1469;
  assign rf_a_tile_v_3_MPORT_45_addr = 8'h32;
  assign rf_a_tile_v_3_MPORT_45_data = rf[rf_a_tile_v_3_MPORT_45_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_2_MPORT_45_en = handshaked & _GEN_1469;
  assign rf_a_tile_v_2_MPORT_45_addr = 8'h36;
  assign rf_a_tile_v_2_MPORT_45_data = rf[rf_a_tile_v_2_MPORT_45_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_1_MPORT_135_en = handshaked & _GEN_1469;
  assign rf_a_tile_v_1_MPORT_135_addr = 8'h3a;
  assign rf_a_tile_v_1_MPORT_135_data = rf[rf_a_tile_v_1_MPORT_135_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_0_MPORT_135_en = handshaked & _GEN_1469;
  assign rf_a_tile_v_0_MPORT_135_addr = 8'h3e;
  assign rf_a_tile_v_0_MPORT_135_data = rf[rf_a_tile_v_0_MPORT_135_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_5_tile_v_3_MPORT_15_en = handshaked & _GEN_1469;
  assign rf_matrix_b_5_tile_v_3_MPORT_15_addr = 8'h61;
  assign rf_matrix_b_5_tile_v_3_MPORT_15_data = rf[rf_matrix_b_5_tile_v_3_MPORT_15_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_5_tile_v_2_MPORT_15_en = handshaked & _GEN_1469;
  assign rf_matrix_b_5_tile_v_2_MPORT_15_addr = 8'h65;
  assign rf_matrix_b_5_tile_v_2_MPORT_15_data = rf[rf_matrix_b_5_tile_v_2_MPORT_15_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_5_tile_v_1_MPORT_15_en = handshaked & _GEN_1469;
  assign rf_matrix_b_5_tile_v_1_MPORT_15_addr = 8'h69;
  assign rf_matrix_b_5_tile_v_1_MPORT_15_data = rf[rf_matrix_b_5_tile_v_1_MPORT_15_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_5_tile_v_0_MPORT_15_en = handshaked & _GEN_1469;
  assign rf_matrix_b_5_tile_v_0_MPORT_15_addr = 8'h6d;
  assign rf_matrix_b_5_tile_v_0_MPORT_15_data = rf[rf_matrix_b_5_tile_v_0_MPORT_15_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_5_tile_v_3_MPORT_15_en = handshaked & _GEN_1469;
  assign rf_matrix_c_5_tile_v_3_MPORT_15_addr = 8'hb1;
  assign rf_matrix_c_5_tile_v_3_MPORT_15_data = rf[rf_matrix_c_5_tile_v_3_MPORT_15_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_5_tile_v_2_MPORT_15_en = handshaked & _GEN_1469;
  assign rf_matrix_c_5_tile_v_2_MPORT_15_addr = 8'hb5;
  assign rf_matrix_c_5_tile_v_2_MPORT_15_data = rf[rf_matrix_c_5_tile_v_2_MPORT_15_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_5_tile_v_1_MPORT_15_en = handshaked & _GEN_1469;
  assign rf_matrix_c_5_tile_v_1_MPORT_15_addr = 8'hb9;
  assign rf_matrix_c_5_tile_v_1_MPORT_15_data = rf[rf_matrix_c_5_tile_v_1_MPORT_15_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_5_tile_v_0_MPORT_15_en = handshaked & _GEN_1469;
  assign rf_matrix_c_5_tile_v_0_MPORT_15_addr = 8'hbd;
  assign rf_matrix_c_5_tile_v_0_MPORT_15_data = rf[rf_matrix_c_5_tile_v_0_MPORT_15_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_1_MPORT_136_en = handshaked & _GEN_1483;
  assign rf_a_tile_v_1_MPORT_136_addr = 8'h32;
  assign rf_a_tile_v_1_MPORT_136_data = rf[rf_a_tile_v_1_MPORT_136_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_0_MPORT_136_en = handshaked & _GEN_1483;
  assign rf_a_tile_v_0_MPORT_136_addr = 8'h36;
  assign rf_a_tile_v_0_MPORT_136_data = rf[rf_a_tile_v_0_MPORT_136_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_5_tile_v_3_MPORT_16_en = handshaked & _GEN_1483;
  assign rf_matrix_b_5_tile_v_3_MPORT_16_addr = 8'h61;
  assign rf_matrix_b_5_tile_v_3_MPORT_16_data = rf[rf_matrix_b_5_tile_v_3_MPORT_16_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_5_tile_v_2_MPORT_16_en = handshaked & _GEN_1483;
  assign rf_matrix_b_5_tile_v_2_MPORT_16_addr = 8'h65;
  assign rf_matrix_b_5_tile_v_2_MPORT_16_data = rf[rf_matrix_b_5_tile_v_2_MPORT_16_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_5_tile_v_1_MPORT_16_en = handshaked & _GEN_1483;
  assign rf_matrix_b_5_tile_v_1_MPORT_16_addr = 8'h69;
  assign rf_matrix_b_5_tile_v_1_MPORT_16_data = rf[rf_matrix_b_5_tile_v_1_MPORT_16_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_5_tile_v_0_MPORT_16_en = handshaked & _GEN_1483;
  assign rf_matrix_b_5_tile_v_0_MPORT_16_addr = 8'h6d;
  assign rf_matrix_b_5_tile_v_0_MPORT_16_data = rf[rf_matrix_b_5_tile_v_0_MPORT_16_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_5_tile_v_3_MPORT_16_en = handshaked & _GEN_1483;
  assign rf_matrix_c_5_tile_v_3_MPORT_16_addr = 8'he2;
  assign rf_matrix_c_5_tile_v_3_MPORT_16_data = rf[rf_matrix_c_5_tile_v_3_MPORT_16_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_5_tile_v_2_MPORT_16_en = handshaked & _GEN_1483;
  assign rf_matrix_c_5_tile_v_2_MPORT_16_addr = 8'he3;
  assign rf_matrix_c_5_tile_v_2_MPORT_16_data = rf[rf_matrix_c_5_tile_v_2_MPORT_16_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_5_tile_v_1_MPORT_16_en = handshaked & _GEN_1483;
  assign rf_matrix_c_5_tile_v_1_MPORT_16_addr = 8'hea;
  assign rf_matrix_c_5_tile_v_1_MPORT_16_data = rf[rf_matrix_c_5_tile_v_1_MPORT_16_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_5_tile_v_0_MPORT_16_en = handshaked & _GEN_1483;
  assign rf_matrix_c_5_tile_v_0_MPORT_16_addr = 8'heb;
  assign rf_matrix_c_5_tile_v_0_MPORT_16_data = rf[rf_matrix_c_5_tile_v_0_MPORT_16_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_1_MPORT_137_en = handshaked & _GEN_1495;
  assign rf_a_tile_v_1_MPORT_137_addr = 8'h3a;
  assign rf_a_tile_v_1_MPORT_137_data = rf[rf_a_tile_v_1_MPORT_137_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_0_MPORT_137_en = handshaked & _GEN_1495;
  assign rf_a_tile_v_0_MPORT_137_addr = 8'h3e;
  assign rf_a_tile_v_0_MPORT_137_data = rf[rf_a_tile_v_0_MPORT_137_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_5_tile_v_3_MPORT_17_en = handshaked & _GEN_1495;
  assign rf_matrix_b_5_tile_v_3_MPORT_17_addr = 8'h61;
  assign rf_matrix_b_5_tile_v_3_MPORT_17_data = rf[rf_matrix_b_5_tile_v_3_MPORT_17_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_5_tile_v_2_MPORT_17_en = handshaked & _GEN_1495;
  assign rf_matrix_b_5_tile_v_2_MPORT_17_addr = 8'h65;
  assign rf_matrix_b_5_tile_v_2_MPORT_17_data = rf[rf_matrix_b_5_tile_v_2_MPORT_17_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_5_tile_v_1_MPORT_17_en = handshaked & _GEN_1495;
  assign rf_matrix_b_5_tile_v_1_MPORT_17_addr = 8'h69;
  assign rf_matrix_b_5_tile_v_1_MPORT_17_data = rf[rf_matrix_b_5_tile_v_1_MPORT_17_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_5_tile_v_0_MPORT_17_en = handshaked & _GEN_1495;
  assign rf_matrix_b_5_tile_v_0_MPORT_17_addr = 8'h6d;
  assign rf_matrix_b_5_tile_v_0_MPORT_17_data = rf[rf_matrix_b_5_tile_v_0_MPORT_17_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_5_tile_v_3_MPORT_17_en = handshaked & _GEN_1495;
  assign rf_matrix_c_5_tile_v_3_MPORT_17_addr = 8'hf2;
  assign rf_matrix_c_5_tile_v_3_MPORT_17_data = rf[rf_matrix_c_5_tile_v_3_MPORT_17_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_5_tile_v_2_MPORT_17_en = handshaked & _GEN_1495;
  assign rf_matrix_c_5_tile_v_2_MPORT_17_addr = 8'hf3;
  assign rf_matrix_c_5_tile_v_2_MPORT_17_data = rf[rf_matrix_c_5_tile_v_2_MPORT_17_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_5_tile_v_1_MPORT_17_en = handshaked & _GEN_1495;
  assign rf_matrix_c_5_tile_v_1_MPORT_17_addr = 8'hfa;
  assign rf_matrix_c_5_tile_v_1_MPORT_17_data = rf[rf_matrix_c_5_tile_v_1_MPORT_17_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_5_tile_v_0_MPORT_17_en = handshaked & _GEN_1495;
  assign rf_matrix_c_5_tile_v_0_MPORT_17_addr = 8'hfb;
  assign rf_matrix_c_5_tile_v_0_MPORT_17_data = rf[rf_matrix_c_5_tile_v_0_MPORT_17_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_1_MPORT_138_en = handshaked & _GEN_1507;
  assign rf_a_tile_v_1_MPORT_138_addr = 8'h33;
  assign rf_a_tile_v_1_MPORT_138_data = rf[rf_a_tile_v_1_MPORT_138_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_0_MPORT_138_en = handshaked & _GEN_1507;
  assign rf_a_tile_v_0_MPORT_138_addr = 8'h37;
  assign rf_a_tile_v_0_MPORT_138_data = rf[rf_a_tile_v_0_MPORT_138_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_5_tile_v_3_MPORT_18_en = handshaked & _GEN_1507;
  assign rf_matrix_b_5_tile_v_3_MPORT_18_addr = 8'h71;
  assign rf_matrix_b_5_tile_v_3_MPORT_18_data = rf[rf_matrix_b_5_tile_v_3_MPORT_18_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_5_tile_v_2_MPORT_18_en = handshaked & _GEN_1507;
  assign rf_matrix_b_5_tile_v_2_MPORT_18_addr = 8'h75;
  assign rf_matrix_b_5_tile_v_2_MPORT_18_data = rf[rf_matrix_b_5_tile_v_2_MPORT_18_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_5_tile_v_1_MPORT_18_en = handshaked & _GEN_1507;
  assign rf_matrix_b_5_tile_v_1_MPORT_18_addr = 8'h79;
  assign rf_matrix_b_5_tile_v_1_MPORT_18_data = rf[rf_matrix_b_5_tile_v_1_MPORT_18_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_5_tile_v_0_MPORT_18_en = handshaked & _GEN_1507;
  assign rf_matrix_b_5_tile_v_0_MPORT_18_addr = 8'h7d;
  assign rf_matrix_b_5_tile_v_0_MPORT_18_data = rf[rf_matrix_b_5_tile_v_0_MPORT_18_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_5_tile_v_3_MPORT_18_en = handshaked & _GEN_1507;
  assign rf_matrix_c_5_tile_v_3_MPORT_18_addr = 8'he0;
  assign rf_matrix_c_5_tile_v_3_MPORT_18_data = rf[rf_matrix_c_5_tile_v_3_MPORT_18_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_5_tile_v_2_MPORT_18_en = handshaked & _GEN_1507;
  assign rf_matrix_c_5_tile_v_2_MPORT_18_addr = 8'he1;
  assign rf_matrix_c_5_tile_v_2_MPORT_18_data = rf[rf_matrix_c_5_tile_v_2_MPORT_18_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_5_tile_v_1_MPORT_18_en = handshaked & _GEN_1507;
  assign rf_matrix_c_5_tile_v_1_MPORT_18_addr = 8'he8;
  assign rf_matrix_c_5_tile_v_1_MPORT_18_data = rf[rf_matrix_c_5_tile_v_1_MPORT_18_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_5_tile_v_0_MPORT_18_en = handshaked & _GEN_1507;
  assign rf_matrix_c_5_tile_v_0_MPORT_18_addr = 8'he9;
  assign rf_matrix_c_5_tile_v_0_MPORT_18_data = rf[rf_matrix_c_5_tile_v_0_MPORT_18_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_3_MPORT_46_en = handshaked & _GEN_1519;
  assign rf_a_tile_v_3_MPORT_46_addr = 8'h33;
  assign rf_a_tile_v_3_MPORT_46_data = rf[rf_a_tile_v_3_MPORT_46_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_2_MPORT_46_en = handshaked & _GEN_1519;
  assign rf_a_tile_v_2_MPORT_46_addr = 8'h37;
  assign rf_a_tile_v_2_MPORT_46_data = rf[rf_a_tile_v_2_MPORT_46_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_1_MPORT_139_en = handshaked & _GEN_1519;
  assign rf_a_tile_v_1_MPORT_139_addr = 8'h3b;
  assign rf_a_tile_v_1_MPORT_139_data = rf[rf_a_tile_v_1_MPORT_139_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_0_MPORT_139_en = handshaked & _GEN_1519;
  assign rf_a_tile_v_0_MPORT_139_addr = 8'h3f;
  assign rf_a_tile_v_0_MPORT_139_data = rf[rf_a_tile_v_0_MPORT_139_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_5_tile_v_3_MPORT_19_en = handshaked & _GEN_1519;
  assign rf_matrix_b_5_tile_v_3_MPORT_19_addr = 8'h71;
  assign rf_matrix_b_5_tile_v_3_MPORT_19_data = rf[rf_matrix_b_5_tile_v_3_MPORT_19_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_5_tile_v_2_MPORT_19_en = handshaked & _GEN_1519;
  assign rf_matrix_b_5_tile_v_2_MPORT_19_addr = 8'h75;
  assign rf_matrix_b_5_tile_v_2_MPORT_19_data = rf[rf_matrix_b_5_tile_v_2_MPORT_19_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_5_tile_v_1_MPORT_19_en = handshaked & _GEN_1519;
  assign rf_matrix_b_5_tile_v_1_MPORT_19_addr = 8'h79;
  assign rf_matrix_b_5_tile_v_1_MPORT_19_data = rf[rf_matrix_b_5_tile_v_1_MPORT_19_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_5_tile_v_0_MPORT_19_en = handshaked & _GEN_1519;
  assign rf_matrix_b_5_tile_v_0_MPORT_19_addr = 8'h7d;
  assign rf_matrix_b_5_tile_v_0_MPORT_19_data = rf[rf_matrix_b_5_tile_v_0_MPORT_19_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_5_tile_v_3_MPORT_19_en = handshaked & _GEN_1519;
  assign rf_matrix_c_5_tile_v_3_MPORT_19_addr = 8'hb0;
  assign rf_matrix_c_5_tile_v_3_MPORT_19_data = rf[rf_matrix_c_5_tile_v_3_MPORT_19_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_5_tile_v_2_MPORT_19_en = handshaked & _GEN_1519;
  assign rf_matrix_c_5_tile_v_2_MPORT_19_addr = 8'hb4;
  assign rf_matrix_c_5_tile_v_2_MPORT_19_data = rf[rf_matrix_c_5_tile_v_2_MPORT_19_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_5_tile_v_1_MPORT_19_en = handshaked & _GEN_1519;
  assign rf_matrix_c_5_tile_v_1_MPORT_19_addr = 8'hb8;
  assign rf_matrix_c_5_tile_v_1_MPORT_19_data = rf[rf_matrix_c_5_tile_v_1_MPORT_19_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_5_tile_v_0_MPORT_19_en = handshaked & _GEN_1519;
  assign rf_matrix_c_5_tile_v_0_MPORT_19_addr = 8'hbc;
  assign rf_matrix_c_5_tile_v_0_MPORT_19_data = rf[rf_matrix_c_5_tile_v_0_MPORT_19_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_1_MPORT_140_en = handshaked & _GEN_1533;
  assign rf_a_tile_v_1_MPORT_140_addr = 8'h3b;
  assign rf_a_tile_v_1_MPORT_140_data = rf[rf_a_tile_v_1_MPORT_140_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_0_MPORT_140_en = handshaked & _GEN_1533;
  assign rf_a_tile_v_0_MPORT_140_addr = 8'h3f;
  assign rf_a_tile_v_0_MPORT_140_data = rf[rf_a_tile_v_0_MPORT_140_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_5_tile_v_3_MPORT_20_en = handshaked & _GEN_1533;
  assign rf_matrix_b_5_tile_v_3_MPORT_20_addr = 8'h71;
  assign rf_matrix_b_5_tile_v_3_MPORT_20_data = rf[rf_matrix_b_5_tile_v_3_MPORT_20_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_5_tile_v_2_MPORT_20_en = handshaked & _GEN_1533;
  assign rf_matrix_b_5_tile_v_2_MPORT_20_addr = 8'h75;
  assign rf_matrix_b_5_tile_v_2_MPORT_20_data = rf[rf_matrix_b_5_tile_v_2_MPORT_20_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_5_tile_v_1_MPORT_20_en = handshaked & _GEN_1533;
  assign rf_matrix_b_5_tile_v_1_MPORT_20_addr = 8'h79;
  assign rf_matrix_b_5_tile_v_1_MPORT_20_data = rf[rf_matrix_b_5_tile_v_1_MPORT_20_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_5_tile_v_0_MPORT_20_en = handshaked & _GEN_1533;
  assign rf_matrix_b_5_tile_v_0_MPORT_20_addr = 8'h7d;
  assign rf_matrix_b_5_tile_v_0_MPORT_20_data = rf[rf_matrix_b_5_tile_v_0_MPORT_20_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_5_tile_v_3_MPORT_20_en = handshaked & _GEN_1533;
  assign rf_matrix_c_5_tile_v_3_MPORT_20_addr = 8'hf0;
  assign rf_matrix_c_5_tile_v_3_MPORT_20_data = rf[rf_matrix_c_5_tile_v_3_MPORT_20_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_5_tile_v_2_MPORT_20_en = handshaked & _GEN_1533;
  assign rf_matrix_c_5_tile_v_2_MPORT_20_addr = 8'hf1;
  assign rf_matrix_c_5_tile_v_2_MPORT_20_data = rf[rf_matrix_c_5_tile_v_2_MPORT_20_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_5_tile_v_1_MPORT_20_en = handshaked & _GEN_1533;
  assign rf_matrix_c_5_tile_v_1_MPORT_20_addr = 8'hf8;
  assign rf_matrix_c_5_tile_v_1_MPORT_20_data = rf[rf_matrix_c_5_tile_v_1_MPORT_20_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_5_tile_v_0_MPORT_20_en = handshaked & _GEN_1533;
  assign rf_matrix_c_5_tile_v_0_MPORT_20_addr = 8'hf9;
  assign rf_matrix_c_5_tile_v_0_MPORT_20_data = rf[rf_matrix_c_5_tile_v_0_MPORT_20_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_3_MPORT_47_en = handshaked & _GEN_1545;
  assign rf_a_tile_v_3_MPORT_47_addr = 8'h33;
  assign rf_a_tile_v_3_MPORT_47_data = rf[rf_a_tile_v_3_MPORT_47_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_2_MPORT_47_en = handshaked & _GEN_1545;
  assign rf_a_tile_v_2_MPORT_47_addr = 8'h37;
  assign rf_a_tile_v_2_MPORT_47_data = rf[rf_a_tile_v_2_MPORT_47_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_1_MPORT_141_en = handshaked & _GEN_1545;
  assign rf_a_tile_v_1_MPORT_141_addr = 8'h3b;
  assign rf_a_tile_v_1_MPORT_141_data = rf[rf_a_tile_v_1_MPORT_141_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_0_MPORT_141_en = handshaked & _GEN_1545;
  assign rf_a_tile_v_0_MPORT_141_addr = 8'h3f;
  assign rf_a_tile_v_0_MPORT_141_data = rf[rf_a_tile_v_0_MPORT_141_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_5_tile_v_3_MPORT_21_en = handshaked & _GEN_1545;
  assign rf_matrix_b_5_tile_v_3_MPORT_21_addr = 8'h71;
  assign rf_matrix_b_5_tile_v_3_MPORT_21_data = rf[rf_matrix_b_5_tile_v_3_MPORT_21_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_5_tile_v_2_MPORT_21_en = handshaked & _GEN_1545;
  assign rf_matrix_b_5_tile_v_2_MPORT_21_addr = 8'h75;
  assign rf_matrix_b_5_tile_v_2_MPORT_21_data = rf[rf_matrix_b_5_tile_v_2_MPORT_21_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_5_tile_v_1_MPORT_21_en = handshaked & _GEN_1545;
  assign rf_matrix_b_5_tile_v_1_MPORT_21_addr = 8'h79;
  assign rf_matrix_b_5_tile_v_1_MPORT_21_data = rf[rf_matrix_b_5_tile_v_1_MPORT_21_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_5_tile_v_0_MPORT_21_en = handshaked & _GEN_1545;
  assign rf_matrix_b_5_tile_v_0_MPORT_21_addr = 8'h7d;
  assign rf_matrix_b_5_tile_v_0_MPORT_21_data = rf[rf_matrix_b_5_tile_v_0_MPORT_21_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_5_tile_v_3_MPORT_21_en = handshaked & _GEN_1545;
  assign rf_matrix_c_5_tile_v_3_MPORT_21_addr = 8'hb1;
  assign rf_matrix_c_5_tile_v_3_MPORT_21_data = rf[rf_matrix_c_5_tile_v_3_MPORT_21_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_5_tile_v_2_MPORT_21_en = handshaked & _GEN_1545;
  assign rf_matrix_c_5_tile_v_2_MPORT_21_addr = 8'hb5;
  assign rf_matrix_c_5_tile_v_2_MPORT_21_data = rf[rf_matrix_c_5_tile_v_2_MPORT_21_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_5_tile_v_1_MPORT_21_en = handshaked & _GEN_1545;
  assign rf_matrix_c_5_tile_v_1_MPORT_21_addr = 8'hb9;
  assign rf_matrix_c_5_tile_v_1_MPORT_21_data = rf[rf_matrix_c_5_tile_v_1_MPORT_21_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_5_tile_v_0_MPORT_21_en = handshaked & _GEN_1545;
  assign rf_matrix_c_5_tile_v_0_MPORT_21_addr = 8'hbd;
  assign rf_matrix_c_5_tile_v_0_MPORT_21_data = rf[rf_matrix_c_5_tile_v_0_MPORT_21_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_1_MPORT_142_en = handshaked & _GEN_1559;
  assign rf_a_tile_v_1_MPORT_142_addr = 8'h33;
  assign rf_a_tile_v_1_MPORT_142_data = rf[rf_a_tile_v_1_MPORT_142_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_0_MPORT_142_en = handshaked & _GEN_1559;
  assign rf_a_tile_v_0_MPORT_142_addr = 8'h37;
  assign rf_a_tile_v_0_MPORT_142_data = rf[rf_a_tile_v_0_MPORT_142_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_5_tile_v_3_MPORT_22_en = handshaked & _GEN_1559;
  assign rf_matrix_b_5_tile_v_3_MPORT_22_addr = 8'h71;
  assign rf_matrix_b_5_tile_v_3_MPORT_22_data = rf[rf_matrix_b_5_tile_v_3_MPORT_22_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_5_tile_v_2_MPORT_22_en = handshaked & _GEN_1559;
  assign rf_matrix_b_5_tile_v_2_MPORT_22_addr = 8'h75;
  assign rf_matrix_b_5_tile_v_2_MPORT_22_data = rf[rf_matrix_b_5_tile_v_2_MPORT_22_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_5_tile_v_1_MPORT_22_en = handshaked & _GEN_1559;
  assign rf_matrix_b_5_tile_v_1_MPORT_22_addr = 8'h79;
  assign rf_matrix_b_5_tile_v_1_MPORT_22_data = rf[rf_matrix_b_5_tile_v_1_MPORT_22_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_5_tile_v_0_MPORT_22_en = handshaked & _GEN_1559;
  assign rf_matrix_b_5_tile_v_0_MPORT_22_addr = 8'h7d;
  assign rf_matrix_b_5_tile_v_0_MPORT_22_data = rf[rf_matrix_b_5_tile_v_0_MPORT_22_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_5_tile_v_3_MPORT_22_en = handshaked & _GEN_1559;
  assign rf_matrix_c_5_tile_v_3_MPORT_22_addr = 8'he2;
  assign rf_matrix_c_5_tile_v_3_MPORT_22_data = rf[rf_matrix_c_5_tile_v_3_MPORT_22_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_5_tile_v_2_MPORT_22_en = handshaked & _GEN_1559;
  assign rf_matrix_c_5_tile_v_2_MPORT_22_addr = 8'he3;
  assign rf_matrix_c_5_tile_v_2_MPORT_22_data = rf[rf_matrix_c_5_tile_v_2_MPORT_22_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_5_tile_v_1_MPORT_22_en = handshaked & _GEN_1559;
  assign rf_matrix_c_5_tile_v_1_MPORT_22_addr = 8'hea;
  assign rf_matrix_c_5_tile_v_1_MPORT_22_data = rf[rf_matrix_c_5_tile_v_1_MPORT_22_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_5_tile_v_0_MPORT_22_en = handshaked & _GEN_1559;
  assign rf_matrix_c_5_tile_v_0_MPORT_22_addr = 8'heb;
  assign rf_matrix_c_5_tile_v_0_MPORT_22_data = rf[rf_matrix_c_5_tile_v_0_MPORT_22_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_1_MPORT_143_en = handshaked & _GEN_1571;
  assign rf_a_tile_v_1_MPORT_143_addr = 8'h3b;
  assign rf_a_tile_v_1_MPORT_143_data = rf[rf_a_tile_v_1_MPORT_143_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_0_MPORT_143_en = handshaked & _GEN_1571;
  assign rf_a_tile_v_0_MPORT_143_addr = 8'h3f;
  assign rf_a_tile_v_0_MPORT_143_data = rf[rf_a_tile_v_0_MPORT_143_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_5_tile_v_3_MPORT_23_en = handshaked & _GEN_1571;
  assign rf_matrix_b_5_tile_v_3_MPORT_23_addr = 8'h71;
  assign rf_matrix_b_5_tile_v_3_MPORT_23_data = rf[rf_matrix_b_5_tile_v_3_MPORT_23_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_5_tile_v_2_MPORT_23_en = handshaked & _GEN_1571;
  assign rf_matrix_b_5_tile_v_2_MPORT_23_addr = 8'h75;
  assign rf_matrix_b_5_tile_v_2_MPORT_23_data = rf[rf_matrix_b_5_tile_v_2_MPORT_23_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_5_tile_v_1_MPORT_23_en = handshaked & _GEN_1571;
  assign rf_matrix_b_5_tile_v_1_MPORT_23_addr = 8'h79;
  assign rf_matrix_b_5_tile_v_1_MPORT_23_data = rf[rf_matrix_b_5_tile_v_1_MPORT_23_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_5_tile_v_0_MPORT_23_en = handshaked & _GEN_1571;
  assign rf_matrix_b_5_tile_v_0_MPORT_23_addr = 8'h7d;
  assign rf_matrix_b_5_tile_v_0_MPORT_23_data = rf[rf_matrix_b_5_tile_v_0_MPORT_23_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_5_tile_v_3_MPORT_23_en = handshaked & _GEN_1571;
  assign rf_matrix_c_5_tile_v_3_MPORT_23_addr = 8'hf2;
  assign rf_matrix_c_5_tile_v_3_MPORT_23_data = rf[rf_matrix_c_5_tile_v_3_MPORT_23_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_5_tile_v_2_MPORT_23_en = handshaked & _GEN_1571;
  assign rf_matrix_c_5_tile_v_2_MPORT_23_addr = 8'hf3;
  assign rf_matrix_c_5_tile_v_2_MPORT_23_data = rf[rf_matrix_c_5_tile_v_2_MPORT_23_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_5_tile_v_1_MPORT_23_en = handshaked & _GEN_1571;
  assign rf_matrix_c_5_tile_v_1_MPORT_23_addr = 8'hfa;
  assign rf_matrix_c_5_tile_v_1_MPORT_23_data = rf[rf_matrix_c_5_tile_v_1_MPORT_23_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_5_tile_v_0_MPORT_23_en = handshaked & _GEN_1571;
  assign rf_matrix_c_5_tile_v_0_MPORT_23_addr = 8'hfb;
  assign rf_matrix_c_5_tile_v_0_MPORT_23_data = rf[rf_matrix_c_5_tile_v_0_MPORT_23_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_1_MPORT_144_en = handshaked & _GEN_1276;
  assign rf_a_tile_v_1_MPORT_144_addr = 8'h10;
  assign rf_a_tile_v_1_MPORT_144_data = rf[rf_a_tile_v_1_MPORT_144_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_0_MPORT_144_en = handshaked & _GEN_1276;
  assign rf_a_tile_v_0_MPORT_144_addr = 8'h14;
  assign rf_a_tile_v_0_MPORT_144_data = rf[rf_a_tile_v_0_MPORT_144_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_6_tile_v_3_MPORT_en = handshaked & _GEN_1276;
  assign rf_matrix_b_6_tile_v_3_MPORT_addr = 8'h43;
  assign rf_matrix_b_6_tile_v_3_MPORT_data = rf[rf_matrix_b_6_tile_v_3_MPORT_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_6_tile_v_2_MPORT_en = handshaked & _GEN_1276;
  assign rf_matrix_b_6_tile_v_2_MPORT_addr = 8'h47;
  assign rf_matrix_b_6_tile_v_2_MPORT_data = rf[rf_matrix_b_6_tile_v_2_MPORT_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_6_tile_v_1_MPORT_en = handshaked & _GEN_1276;
  assign rf_matrix_b_6_tile_v_1_MPORT_addr = 8'h4b;
  assign rf_matrix_b_6_tile_v_1_MPORT_data = rf[rf_matrix_b_6_tile_v_1_MPORT_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_6_tile_v_0_MPORT_en = handshaked & _GEN_1276;
  assign rf_matrix_b_6_tile_v_0_MPORT_addr = 8'h4f;
  assign rf_matrix_b_6_tile_v_0_MPORT_data = rf[rf_matrix_b_6_tile_v_0_MPORT_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_6_tile_v_3_MPORT_en = handshaked & _GEN_1276;
  assign rf_matrix_c_6_tile_v_3_MPORT_addr = 8'ha4;
  assign rf_matrix_c_6_tile_v_3_MPORT_data = rf[rf_matrix_c_6_tile_v_3_MPORT_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_6_tile_v_2_MPORT_en = handshaked & _GEN_1276;
  assign rf_matrix_c_6_tile_v_2_MPORT_addr = 8'ha5;
  assign rf_matrix_c_6_tile_v_2_MPORT_data = rf[rf_matrix_c_6_tile_v_2_MPORT_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_6_tile_v_1_MPORT_en = handshaked & _GEN_1276;
  assign rf_matrix_c_6_tile_v_1_MPORT_addr = 8'hac;
  assign rf_matrix_c_6_tile_v_1_MPORT_data = rf[rf_matrix_c_6_tile_v_1_MPORT_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_6_tile_v_0_MPORT_en = handshaked & _GEN_1276;
  assign rf_matrix_c_6_tile_v_0_MPORT_addr = 8'had;
  assign rf_matrix_c_6_tile_v_0_MPORT_data = rf[rf_matrix_c_6_tile_v_0_MPORT_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_3_MPORT_48_en = handshaked & _GEN_1291;
  assign rf_a_tile_v_3_MPORT_48_addr = 8'h10;
  assign rf_a_tile_v_3_MPORT_48_data = rf[rf_a_tile_v_3_MPORT_48_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_2_MPORT_48_en = handshaked & _GEN_1291;
  assign rf_a_tile_v_2_MPORT_48_addr = 8'h14;
  assign rf_a_tile_v_2_MPORT_48_data = rf[rf_a_tile_v_2_MPORT_48_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_1_MPORT_145_en = handshaked & _GEN_1291;
  assign rf_a_tile_v_1_MPORT_145_addr = 8'h18;
  assign rf_a_tile_v_1_MPORT_145_data = rf[rf_a_tile_v_1_MPORT_145_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_0_MPORT_145_en = handshaked & _GEN_1291;
  assign rf_a_tile_v_0_MPORT_145_addr = 8'h1c;
  assign rf_a_tile_v_0_MPORT_145_data = rf[rf_a_tile_v_0_MPORT_145_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_6_tile_v_3_MPORT_1_en = handshaked & _GEN_1291;
  assign rf_matrix_b_6_tile_v_3_MPORT_1_addr = 8'h43;
  assign rf_matrix_b_6_tile_v_3_MPORT_1_data = rf[rf_matrix_b_6_tile_v_3_MPORT_1_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_6_tile_v_2_MPORT_1_en = handshaked & _GEN_1291;
  assign rf_matrix_b_6_tile_v_2_MPORT_1_addr = 8'h47;
  assign rf_matrix_b_6_tile_v_2_MPORT_1_data = rf[rf_matrix_b_6_tile_v_2_MPORT_1_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_6_tile_v_1_MPORT_1_en = handshaked & _GEN_1291;
  assign rf_matrix_b_6_tile_v_1_MPORT_1_addr = 8'h4b;
  assign rf_matrix_b_6_tile_v_1_MPORT_1_data = rf[rf_matrix_b_6_tile_v_1_MPORT_1_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_6_tile_v_0_MPORT_1_en = handshaked & _GEN_1291;
  assign rf_matrix_b_6_tile_v_0_MPORT_1_addr = 8'h4f;
  assign rf_matrix_b_6_tile_v_0_MPORT_1_data = rf[rf_matrix_b_6_tile_v_0_MPORT_1_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_6_tile_v_3_MPORT_1_en = handshaked & _GEN_1291;
  assign rf_matrix_c_6_tile_v_3_MPORT_1_addr = 8'h92;
  assign rf_matrix_c_6_tile_v_3_MPORT_1_data = rf[rf_matrix_c_6_tile_v_3_MPORT_1_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_6_tile_v_2_MPORT_1_en = handshaked & _GEN_1291;
  assign rf_matrix_c_6_tile_v_2_MPORT_1_addr = 8'h96;
  assign rf_matrix_c_6_tile_v_2_MPORT_1_data = rf[rf_matrix_c_6_tile_v_2_MPORT_1_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_6_tile_v_1_MPORT_1_en = handshaked & _GEN_1291;
  assign rf_matrix_c_6_tile_v_1_MPORT_1_addr = 8'h9a;
  assign rf_matrix_c_6_tile_v_1_MPORT_1_data = rf[rf_matrix_c_6_tile_v_1_MPORT_1_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_6_tile_v_0_MPORT_1_en = handshaked & _GEN_1291;
  assign rf_matrix_c_6_tile_v_0_MPORT_1_addr = 8'h9e;
  assign rf_matrix_c_6_tile_v_0_MPORT_1_data = rf[rf_matrix_c_6_tile_v_0_MPORT_1_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_1_MPORT_146_en = handshaked & _GEN_1305;
  assign rf_a_tile_v_1_MPORT_146_addr = 8'h18;
  assign rf_a_tile_v_1_MPORT_146_data = rf[rf_a_tile_v_1_MPORT_146_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_0_MPORT_146_en = handshaked & _GEN_1305;
  assign rf_a_tile_v_0_MPORT_146_addr = 8'h1c;
  assign rf_a_tile_v_0_MPORT_146_data = rf[rf_a_tile_v_0_MPORT_146_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_6_tile_v_3_MPORT_2_en = handshaked & _GEN_1305;
  assign rf_matrix_b_6_tile_v_3_MPORT_2_addr = 8'h43;
  assign rf_matrix_b_6_tile_v_3_MPORT_2_data = rf[rf_matrix_b_6_tile_v_3_MPORT_2_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_6_tile_v_2_MPORT_2_en = handshaked & _GEN_1305;
  assign rf_matrix_b_6_tile_v_2_MPORT_2_addr = 8'h47;
  assign rf_matrix_b_6_tile_v_2_MPORT_2_data = rf[rf_matrix_b_6_tile_v_2_MPORT_2_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_6_tile_v_1_MPORT_2_en = handshaked & _GEN_1305;
  assign rf_matrix_b_6_tile_v_1_MPORT_2_addr = 8'h4b;
  assign rf_matrix_b_6_tile_v_1_MPORT_2_data = rf[rf_matrix_b_6_tile_v_1_MPORT_2_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_6_tile_v_0_MPORT_2_en = handshaked & _GEN_1305;
  assign rf_matrix_b_6_tile_v_0_MPORT_2_addr = 8'h4f;
  assign rf_matrix_b_6_tile_v_0_MPORT_2_data = rf[rf_matrix_b_6_tile_v_0_MPORT_2_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_6_tile_v_3_MPORT_2_en = handshaked & _GEN_1305;
  assign rf_matrix_c_6_tile_v_3_MPORT_2_addr = 8'hb4;
  assign rf_matrix_c_6_tile_v_3_MPORT_2_data = rf[rf_matrix_c_6_tile_v_3_MPORT_2_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_6_tile_v_2_MPORT_2_en = handshaked & _GEN_1305;
  assign rf_matrix_c_6_tile_v_2_MPORT_2_addr = 8'hb5;
  assign rf_matrix_c_6_tile_v_2_MPORT_2_data = rf[rf_matrix_c_6_tile_v_2_MPORT_2_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_6_tile_v_1_MPORT_2_en = handshaked & _GEN_1305;
  assign rf_matrix_c_6_tile_v_1_MPORT_2_addr = 8'hbc;
  assign rf_matrix_c_6_tile_v_1_MPORT_2_data = rf[rf_matrix_c_6_tile_v_1_MPORT_2_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_6_tile_v_0_MPORT_2_en = handshaked & _GEN_1305;
  assign rf_matrix_c_6_tile_v_0_MPORT_2_addr = 8'hbd;
  assign rf_matrix_c_6_tile_v_0_MPORT_2_data = rf[rf_matrix_c_6_tile_v_0_MPORT_2_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_3_MPORT_49_en = handshaked & _GEN_1317;
  assign rf_a_tile_v_3_MPORT_49_addr = 8'h10;
  assign rf_a_tile_v_3_MPORT_49_data = rf[rf_a_tile_v_3_MPORT_49_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_2_MPORT_49_en = handshaked & _GEN_1317;
  assign rf_a_tile_v_2_MPORT_49_addr = 8'h14;
  assign rf_a_tile_v_2_MPORT_49_data = rf[rf_a_tile_v_2_MPORT_49_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_1_MPORT_147_en = handshaked & _GEN_1317;
  assign rf_a_tile_v_1_MPORT_147_addr = 8'h18;
  assign rf_a_tile_v_1_MPORT_147_data = rf[rf_a_tile_v_1_MPORT_147_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_0_MPORT_147_en = handshaked & _GEN_1317;
  assign rf_a_tile_v_0_MPORT_147_addr = 8'h1c;
  assign rf_a_tile_v_0_MPORT_147_data = rf[rf_a_tile_v_0_MPORT_147_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_6_tile_v_3_MPORT_3_en = handshaked & _GEN_1317;
  assign rf_matrix_b_6_tile_v_3_MPORT_3_addr = 8'h43;
  assign rf_matrix_b_6_tile_v_3_MPORT_3_data = rf[rf_matrix_b_6_tile_v_3_MPORT_3_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_6_tile_v_2_MPORT_3_en = handshaked & _GEN_1317;
  assign rf_matrix_b_6_tile_v_2_MPORT_3_addr = 8'h47;
  assign rf_matrix_b_6_tile_v_2_MPORT_3_data = rf[rf_matrix_b_6_tile_v_2_MPORT_3_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_6_tile_v_1_MPORT_3_en = handshaked & _GEN_1317;
  assign rf_matrix_b_6_tile_v_1_MPORT_3_addr = 8'h4b;
  assign rf_matrix_b_6_tile_v_1_MPORT_3_data = rf[rf_matrix_b_6_tile_v_1_MPORT_3_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_6_tile_v_0_MPORT_3_en = handshaked & _GEN_1317;
  assign rf_matrix_b_6_tile_v_0_MPORT_3_addr = 8'h4f;
  assign rf_matrix_b_6_tile_v_0_MPORT_3_data = rf[rf_matrix_b_6_tile_v_0_MPORT_3_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_6_tile_v_3_MPORT_3_en = handshaked & _GEN_1317;
  assign rf_matrix_c_6_tile_v_3_MPORT_3_addr = 8'h93;
  assign rf_matrix_c_6_tile_v_3_MPORT_3_data = rf[rf_matrix_c_6_tile_v_3_MPORT_3_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_6_tile_v_2_MPORT_3_en = handshaked & _GEN_1317;
  assign rf_matrix_c_6_tile_v_2_MPORT_3_addr = 8'h97;
  assign rf_matrix_c_6_tile_v_2_MPORT_3_data = rf[rf_matrix_c_6_tile_v_2_MPORT_3_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_6_tile_v_1_MPORT_3_en = handshaked & _GEN_1317;
  assign rf_matrix_c_6_tile_v_1_MPORT_3_addr = 8'h9b;
  assign rf_matrix_c_6_tile_v_1_MPORT_3_data = rf[rf_matrix_c_6_tile_v_1_MPORT_3_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_6_tile_v_0_MPORT_3_en = handshaked & _GEN_1317;
  assign rf_matrix_c_6_tile_v_0_MPORT_3_addr = 8'h9f;
  assign rf_matrix_c_6_tile_v_0_MPORT_3_data = rf[rf_matrix_c_6_tile_v_0_MPORT_3_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_1_MPORT_148_en = handshaked & _GEN_1331;
  assign rf_a_tile_v_1_MPORT_148_addr = 8'h10;
  assign rf_a_tile_v_1_MPORT_148_data = rf[rf_a_tile_v_1_MPORT_148_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_0_MPORT_148_en = handshaked & _GEN_1331;
  assign rf_a_tile_v_0_MPORT_148_addr = 8'h14;
  assign rf_a_tile_v_0_MPORT_148_data = rf[rf_a_tile_v_0_MPORT_148_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_6_tile_v_3_MPORT_4_en = handshaked & _GEN_1331;
  assign rf_matrix_b_6_tile_v_3_MPORT_4_addr = 8'h43;
  assign rf_matrix_b_6_tile_v_3_MPORT_4_data = rf[rf_matrix_b_6_tile_v_3_MPORT_4_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_6_tile_v_2_MPORT_4_en = handshaked & _GEN_1331;
  assign rf_matrix_b_6_tile_v_2_MPORT_4_addr = 8'h47;
  assign rf_matrix_b_6_tile_v_2_MPORT_4_data = rf[rf_matrix_b_6_tile_v_2_MPORT_4_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_6_tile_v_1_MPORT_4_en = handshaked & _GEN_1331;
  assign rf_matrix_b_6_tile_v_1_MPORT_4_addr = 8'h4b;
  assign rf_matrix_b_6_tile_v_1_MPORT_4_data = rf[rf_matrix_b_6_tile_v_1_MPORT_4_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_6_tile_v_0_MPORT_4_en = handshaked & _GEN_1331;
  assign rf_matrix_b_6_tile_v_0_MPORT_4_addr = 8'h4f;
  assign rf_matrix_b_6_tile_v_0_MPORT_4_data = rf[rf_matrix_b_6_tile_v_0_MPORT_4_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_6_tile_v_3_MPORT_4_en = handshaked & _GEN_1331;
  assign rf_matrix_c_6_tile_v_3_MPORT_4_addr = 8'ha6;
  assign rf_matrix_c_6_tile_v_3_MPORT_4_data = rf[rf_matrix_c_6_tile_v_3_MPORT_4_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_6_tile_v_2_MPORT_4_en = handshaked & _GEN_1331;
  assign rf_matrix_c_6_tile_v_2_MPORT_4_addr = 8'ha7;
  assign rf_matrix_c_6_tile_v_2_MPORT_4_data = rf[rf_matrix_c_6_tile_v_2_MPORT_4_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_6_tile_v_1_MPORT_4_en = handshaked & _GEN_1331;
  assign rf_matrix_c_6_tile_v_1_MPORT_4_addr = 8'hae;
  assign rf_matrix_c_6_tile_v_1_MPORT_4_data = rf[rf_matrix_c_6_tile_v_1_MPORT_4_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_6_tile_v_0_MPORT_4_en = handshaked & _GEN_1331;
  assign rf_matrix_c_6_tile_v_0_MPORT_4_addr = 8'haf;
  assign rf_matrix_c_6_tile_v_0_MPORT_4_data = rf[rf_matrix_c_6_tile_v_0_MPORT_4_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_1_MPORT_149_en = handshaked & _GEN_1343;
  assign rf_a_tile_v_1_MPORT_149_addr = 8'h18;
  assign rf_a_tile_v_1_MPORT_149_data = rf[rf_a_tile_v_1_MPORT_149_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_0_MPORT_149_en = handshaked & _GEN_1343;
  assign rf_a_tile_v_0_MPORT_149_addr = 8'h1c;
  assign rf_a_tile_v_0_MPORT_149_data = rf[rf_a_tile_v_0_MPORT_149_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_6_tile_v_3_MPORT_5_en = handshaked & _GEN_1343;
  assign rf_matrix_b_6_tile_v_3_MPORT_5_addr = 8'h43;
  assign rf_matrix_b_6_tile_v_3_MPORT_5_data = rf[rf_matrix_b_6_tile_v_3_MPORT_5_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_6_tile_v_2_MPORT_5_en = handshaked & _GEN_1343;
  assign rf_matrix_b_6_tile_v_2_MPORT_5_addr = 8'h47;
  assign rf_matrix_b_6_tile_v_2_MPORT_5_data = rf[rf_matrix_b_6_tile_v_2_MPORT_5_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_6_tile_v_1_MPORT_5_en = handshaked & _GEN_1343;
  assign rf_matrix_b_6_tile_v_1_MPORT_5_addr = 8'h4b;
  assign rf_matrix_b_6_tile_v_1_MPORT_5_data = rf[rf_matrix_b_6_tile_v_1_MPORT_5_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_6_tile_v_0_MPORT_5_en = handshaked & _GEN_1343;
  assign rf_matrix_b_6_tile_v_0_MPORT_5_addr = 8'h4f;
  assign rf_matrix_b_6_tile_v_0_MPORT_5_data = rf[rf_matrix_b_6_tile_v_0_MPORT_5_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_6_tile_v_3_MPORT_5_en = handshaked & _GEN_1343;
  assign rf_matrix_c_6_tile_v_3_MPORT_5_addr = 8'hb6;
  assign rf_matrix_c_6_tile_v_3_MPORT_5_data = rf[rf_matrix_c_6_tile_v_3_MPORT_5_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_6_tile_v_2_MPORT_5_en = handshaked & _GEN_1343;
  assign rf_matrix_c_6_tile_v_2_MPORT_5_addr = 8'hb7;
  assign rf_matrix_c_6_tile_v_2_MPORT_5_data = rf[rf_matrix_c_6_tile_v_2_MPORT_5_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_6_tile_v_1_MPORT_5_en = handshaked & _GEN_1343;
  assign rf_matrix_c_6_tile_v_1_MPORT_5_addr = 8'hbe;
  assign rf_matrix_c_6_tile_v_1_MPORT_5_data = rf[rf_matrix_c_6_tile_v_1_MPORT_5_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_6_tile_v_0_MPORT_5_en = handshaked & _GEN_1343;
  assign rf_matrix_c_6_tile_v_0_MPORT_5_addr = 8'hbf;
  assign rf_matrix_c_6_tile_v_0_MPORT_5_data = rf[rf_matrix_c_6_tile_v_0_MPORT_5_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_1_MPORT_150_en = handshaked & _GEN_1355;
  assign rf_a_tile_v_1_MPORT_150_addr = 8'h11;
  assign rf_a_tile_v_1_MPORT_150_data = rf[rf_a_tile_v_1_MPORT_150_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_0_MPORT_150_en = handshaked & _GEN_1355;
  assign rf_a_tile_v_0_MPORT_150_addr = 8'h15;
  assign rf_a_tile_v_0_MPORT_150_data = rf[rf_a_tile_v_0_MPORT_150_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_6_tile_v_3_MPORT_6_en = handshaked & _GEN_1355;
  assign rf_matrix_b_6_tile_v_3_MPORT_6_addr = 8'h53;
  assign rf_matrix_b_6_tile_v_3_MPORT_6_data = rf[rf_matrix_b_6_tile_v_3_MPORT_6_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_6_tile_v_2_MPORT_6_en = handshaked & _GEN_1355;
  assign rf_matrix_b_6_tile_v_2_MPORT_6_addr = 8'h57;
  assign rf_matrix_b_6_tile_v_2_MPORT_6_data = rf[rf_matrix_b_6_tile_v_2_MPORT_6_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_6_tile_v_1_MPORT_6_en = handshaked & _GEN_1355;
  assign rf_matrix_b_6_tile_v_1_MPORT_6_addr = 8'h5b;
  assign rf_matrix_b_6_tile_v_1_MPORT_6_data = rf[rf_matrix_b_6_tile_v_1_MPORT_6_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_6_tile_v_0_MPORT_6_en = handshaked & _GEN_1355;
  assign rf_matrix_b_6_tile_v_0_MPORT_6_addr = 8'h5f;
  assign rf_matrix_b_6_tile_v_0_MPORT_6_data = rf[rf_matrix_b_6_tile_v_0_MPORT_6_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_6_tile_v_3_MPORT_6_en = handshaked & _GEN_1355;
  assign rf_matrix_c_6_tile_v_3_MPORT_6_addr = 8'ha4;
  assign rf_matrix_c_6_tile_v_3_MPORT_6_data = rf[rf_matrix_c_6_tile_v_3_MPORT_6_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_6_tile_v_2_MPORT_6_en = handshaked & _GEN_1355;
  assign rf_matrix_c_6_tile_v_2_MPORT_6_addr = 8'ha5;
  assign rf_matrix_c_6_tile_v_2_MPORT_6_data = rf[rf_matrix_c_6_tile_v_2_MPORT_6_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_6_tile_v_1_MPORT_6_en = handshaked & _GEN_1355;
  assign rf_matrix_c_6_tile_v_1_MPORT_6_addr = 8'hac;
  assign rf_matrix_c_6_tile_v_1_MPORT_6_data = rf[rf_matrix_c_6_tile_v_1_MPORT_6_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_6_tile_v_0_MPORT_6_en = handshaked & _GEN_1355;
  assign rf_matrix_c_6_tile_v_0_MPORT_6_addr = 8'had;
  assign rf_matrix_c_6_tile_v_0_MPORT_6_data = rf[rf_matrix_c_6_tile_v_0_MPORT_6_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_3_MPORT_50_en = handshaked & _GEN_1367;
  assign rf_a_tile_v_3_MPORT_50_addr = 8'h11;
  assign rf_a_tile_v_3_MPORT_50_data = rf[rf_a_tile_v_3_MPORT_50_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_2_MPORT_50_en = handshaked & _GEN_1367;
  assign rf_a_tile_v_2_MPORT_50_addr = 8'h15;
  assign rf_a_tile_v_2_MPORT_50_data = rf[rf_a_tile_v_2_MPORT_50_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_1_MPORT_151_en = handshaked & _GEN_1367;
  assign rf_a_tile_v_1_MPORT_151_addr = 8'h19;
  assign rf_a_tile_v_1_MPORT_151_data = rf[rf_a_tile_v_1_MPORT_151_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_0_MPORT_151_en = handshaked & _GEN_1367;
  assign rf_a_tile_v_0_MPORT_151_addr = 8'h1d;
  assign rf_a_tile_v_0_MPORT_151_data = rf[rf_a_tile_v_0_MPORT_151_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_6_tile_v_3_MPORT_7_en = handshaked & _GEN_1367;
  assign rf_matrix_b_6_tile_v_3_MPORT_7_addr = 8'h53;
  assign rf_matrix_b_6_tile_v_3_MPORT_7_data = rf[rf_matrix_b_6_tile_v_3_MPORT_7_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_6_tile_v_2_MPORT_7_en = handshaked & _GEN_1367;
  assign rf_matrix_b_6_tile_v_2_MPORT_7_addr = 8'h57;
  assign rf_matrix_b_6_tile_v_2_MPORT_7_data = rf[rf_matrix_b_6_tile_v_2_MPORT_7_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_6_tile_v_1_MPORT_7_en = handshaked & _GEN_1367;
  assign rf_matrix_b_6_tile_v_1_MPORT_7_addr = 8'h5b;
  assign rf_matrix_b_6_tile_v_1_MPORT_7_data = rf[rf_matrix_b_6_tile_v_1_MPORT_7_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_6_tile_v_0_MPORT_7_en = handshaked & _GEN_1367;
  assign rf_matrix_b_6_tile_v_0_MPORT_7_addr = 8'h5f;
  assign rf_matrix_b_6_tile_v_0_MPORT_7_data = rf[rf_matrix_b_6_tile_v_0_MPORT_7_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_6_tile_v_3_MPORT_7_en = handshaked & _GEN_1367;
  assign rf_matrix_c_6_tile_v_3_MPORT_7_addr = 8'h92;
  assign rf_matrix_c_6_tile_v_3_MPORT_7_data = rf[rf_matrix_c_6_tile_v_3_MPORT_7_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_6_tile_v_2_MPORT_7_en = handshaked & _GEN_1367;
  assign rf_matrix_c_6_tile_v_2_MPORT_7_addr = 8'h96;
  assign rf_matrix_c_6_tile_v_2_MPORT_7_data = rf[rf_matrix_c_6_tile_v_2_MPORT_7_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_6_tile_v_1_MPORT_7_en = handshaked & _GEN_1367;
  assign rf_matrix_c_6_tile_v_1_MPORT_7_addr = 8'h9a;
  assign rf_matrix_c_6_tile_v_1_MPORT_7_data = rf[rf_matrix_c_6_tile_v_1_MPORT_7_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_6_tile_v_0_MPORT_7_en = handshaked & _GEN_1367;
  assign rf_matrix_c_6_tile_v_0_MPORT_7_addr = 8'h9e;
  assign rf_matrix_c_6_tile_v_0_MPORT_7_data = rf[rf_matrix_c_6_tile_v_0_MPORT_7_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_1_MPORT_152_en = handshaked & _GEN_1381;
  assign rf_a_tile_v_1_MPORT_152_addr = 8'h19;
  assign rf_a_tile_v_1_MPORT_152_data = rf[rf_a_tile_v_1_MPORT_152_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_0_MPORT_152_en = handshaked & _GEN_1381;
  assign rf_a_tile_v_0_MPORT_152_addr = 8'h1d;
  assign rf_a_tile_v_0_MPORT_152_data = rf[rf_a_tile_v_0_MPORT_152_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_6_tile_v_3_MPORT_8_en = handshaked & _GEN_1381;
  assign rf_matrix_b_6_tile_v_3_MPORT_8_addr = 8'h53;
  assign rf_matrix_b_6_tile_v_3_MPORT_8_data = rf[rf_matrix_b_6_tile_v_3_MPORT_8_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_6_tile_v_2_MPORT_8_en = handshaked & _GEN_1381;
  assign rf_matrix_b_6_tile_v_2_MPORT_8_addr = 8'h57;
  assign rf_matrix_b_6_tile_v_2_MPORT_8_data = rf[rf_matrix_b_6_tile_v_2_MPORT_8_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_6_tile_v_1_MPORT_8_en = handshaked & _GEN_1381;
  assign rf_matrix_b_6_tile_v_1_MPORT_8_addr = 8'h5b;
  assign rf_matrix_b_6_tile_v_1_MPORT_8_data = rf[rf_matrix_b_6_tile_v_1_MPORT_8_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_6_tile_v_0_MPORT_8_en = handshaked & _GEN_1381;
  assign rf_matrix_b_6_tile_v_0_MPORT_8_addr = 8'h5f;
  assign rf_matrix_b_6_tile_v_0_MPORT_8_data = rf[rf_matrix_b_6_tile_v_0_MPORT_8_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_6_tile_v_3_MPORT_8_en = handshaked & _GEN_1381;
  assign rf_matrix_c_6_tile_v_3_MPORT_8_addr = 8'hb4;
  assign rf_matrix_c_6_tile_v_3_MPORT_8_data = rf[rf_matrix_c_6_tile_v_3_MPORT_8_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_6_tile_v_2_MPORT_8_en = handshaked & _GEN_1381;
  assign rf_matrix_c_6_tile_v_2_MPORT_8_addr = 8'hb5;
  assign rf_matrix_c_6_tile_v_2_MPORT_8_data = rf[rf_matrix_c_6_tile_v_2_MPORT_8_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_6_tile_v_1_MPORT_8_en = handshaked & _GEN_1381;
  assign rf_matrix_c_6_tile_v_1_MPORT_8_addr = 8'hbc;
  assign rf_matrix_c_6_tile_v_1_MPORT_8_data = rf[rf_matrix_c_6_tile_v_1_MPORT_8_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_6_tile_v_0_MPORT_8_en = handshaked & _GEN_1381;
  assign rf_matrix_c_6_tile_v_0_MPORT_8_addr = 8'hbd;
  assign rf_matrix_c_6_tile_v_0_MPORT_8_data = rf[rf_matrix_c_6_tile_v_0_MPORT_8_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_3_MPORT_51_en = handshaked & _GEN_1393;
  assign rf_a_tile_v_3_MPORT_51_addr = 8'h11;
  assign rf_a_tile_v_3_MPORT_51_data = rf[rf_a_tile_v_3_MPORT_51_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_2_MPORT_51_en = handshaked & _GEN_1393;
  assign rf_a_tile_v_2_MPORT_51_addr = 8'h15;
  assign rf_a_tile_v_2_MPORT_51_data = rf[rf_a_tile_v_2_MPORT_51_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_1_MPORT_153_en = handshaked & _GEN_1393;
  assign rf_a_tile_v_1_MPORT_153_addr = 8'h19;
  assign rf_a_tile_v_1_MPORT_153_data = rf[rf_a_tile_v_1_MPORT_153_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_0_MPORT_153_en = handshaked & _GEN_1393;
  assign rf_a_tile_v_0_MPORT_153_addr = 8'h1d;
  assign rf_a_tile_v_0_MPORT_153_data = rf[rf_a_tile_v_0_MPORT_153_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_6_tile_v_3_MPORT_9_en = handshaked & _GEN_1393;
  assign rf_matrix_b_6_tile_v_3_MPORT_9_addr = 8'h53;
  assign rf_matrix_b_6_tile_v_3_MPORT_9_data = rf[rf_matrix_b_6_tile_v_3_MPORT_9_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_6_tile_v_2_MPORT_9_en = handshaked & _GEN_1393;
  assign rf_matrix_b_6_tile_v_2_MPORT_9_addr = 8'h57;
  assign rf_matrix_b_6_tile_v_2_MPORT_9_data = rf[rf_matrix_b_6_tile_v_2_MPORT_9_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_6_tile_v_1_MPORT_9_en = handshaked & _GEN_1393;
  assign rf_matrix_b_6_tile_v_1_MPORT_9_addr = 8'h5b;
  assign rf_matrix_b_6_tile_v_1_MPORT_9_data = rf[rf_matrix_b_6_tile_v_1_MPORT_9_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_6_tile_v_0_MPORT_9_en = handshaked & _GEN_1393;
  assign rf_matrix_b_6_tile_v_0_MPORT_9_addr = 8'h5f;
  assign rf_matrix_b_6_tile_v_0_MPORT_9_data = rf[rf_matrix_b_6_tile_v_0_MPORT_9_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_6_tile_v_3_MPORT_9_en = handshaked & _GEN_1393;
  assign rf_matrix_c_6_tile_v_3_MPORT_9_addr = 8'h93;
  assign rf_matrix_c_6_tile_v_3_MPORT_9_data = rf[rf_matrix_c_6_tile_v_3_MPORT_9_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_6_tile_v_2_MPORT_9_en = handshaked & _GEN_1393;
  assign rf_matrix_c_6_tile_v_2_MPORT_9_addr = 8'h97;
  assign rf_matrix_c_6_tile_v_2_MPORT_9_data = rf[rf_matrix_c_6_tile_v_2_MPORT_9_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_6_tile_v_1_MPORT_9_en = handshaked & _GEN_1393;
  assign rf_matrix_c_6_tile_v_1_MPORT_9_addr = 8'h9b;
  assign rf_matrix_c_6_tile_v_1_MPORT_9_data = rf[rf_matrix_c_6_tile_v_1_MPORT_9_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_6_tile_v_0_MPORT_9_en = handshaked & _GEN_1393;
  assign rf_matrix_c_6_tile_v_0_MPORT_9_addr = 8'h9f;
  assign rf_matrix_c_6_tile_v_0_MPORT_9_data = rf[rf_matrix_c_6_tile_v_0_MPORT_9_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_1_MPORT_154_en = handshaked & _GEN_1407;
  assign rf_a_tile_v_1_MPORT_154_addr = 8'h11;
  assign rf_a_tile_v_1_MPORT_154_data = rf[rf_a_tile_v_1_MPORT_154_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_0_MPORT_154_en = handshaked & _GEN_1407;
  assign rf_a_tile_v_0_MPORT_154_addr = 8'h15;
  assign rf_a_tile_v_0_MPORT_154_data = rf[rf_a_tile_v_0_MPORT_154_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_6_tile_v_3_MPORT_10_en = handshaked & _GEN_1407;
  assign rf_matrix_b_6_tile_v_3_MPORT_10_addr = 8'h53;
  assign rf_matrix_b_6_tile_v_3_MPORT_10_data = rf[rf_matrix_b_6_tile_v_3_MPORT_10_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_6_tile_v_2_MPORT_10_en = handshaked & _GEN_1407;
  assign rf_matrix_b_6_tile_v_2_MPORT_10_addr = 8'h57;
  assign rf_matrix_b_6_tile_v_2_MPORT_10_data = rf[rf_matrix_b_6_tile_v_2_MPORT_10_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_6_tile_v_1_MPORT_10_en = handshaked & _GEN_1407;
  assign rf_matrix_b_6_tile_v_1_MPORT_10_addr = 8'h5b;
  assign rf_matrix_b_6_tile_v_1_MPORT_10_data = rf[rf_matrix_b_6_tile_v_1_MPORT_10_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_6_tile_v_0_MPORT_10_en = handshaked & _GEN_1407;
  assign rf_matrix_b_6_tile_v_0_MPORT_10_addr = 8'h5f;
  assign rf_matrix_b_6_tile_v_0_MPORT_10_data = rf[rf_matrix_b_6_tile_v_0_MPORT_10_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_6_tile_v_3_MPORT_10_en = handshaked & _GEN_1407;
  assign rf_matrix_c_6_tile_v_3_MPORT_10_addr = 8'ha6;
  assign rf_matrix_c_6_tile_v_3_MPORT_10_data = rf[rf_matrix_c_6_tile_v_3_MPORT_10_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_6_tile_v_2_MPORT_10_en = handshaked & _GEN_1407;
  assign rf_matrix_c_6_tile_v_2_MPORT_10_addr = 8'ha7;
  assign rf_matrix_c_6_tile_v_2_MPORT_10_data = rf[rf_matrix_c_6_tile_v_2_MPORT_10_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_6_tile_v_1_MPORT_10_en = handshaked & _GEN_1407;
  assign rf_matrix_c_6_tile_v_1_MPORT_10_addr = 8'hae;
  assign rf_matrix_c_6_tile_v_1_MPORT_10_data = rf[rf_matrix_c_6_tile_v_1_MPORT_10_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_6_tile_v_0_MPORT_10_en = handshaked & _GEN_1407;
  assign rf_matrix_c_6_tile_v_0_MPORT_10_addr = 8'haf;
  assign rf_matrix_c_6_tile_v_0_MPORT_10_data = rf[rf_matrix_c_6_tile_v_0_MPORT_10_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_1_MPORT_155_en = handshaked & _GEN_1419;
  assign rf_a_tile_v_1_MPORT_155_addr = 8'h19;
  assign rf_a_tile_v_1_MPORT_155_data = rf[rf_a_tile_v_1_MPORT_155_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_0_MPORT_155_en = handshaked & _GEN_1419;
  assign rf_a_tile_v_0_MPORT_155_addr = 8'h1d;
  assign rf_a_tile_v_0_MPORT_155_data = rf[rf_a_tile_v_0_MPORT_155_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_6_tile_v_3_MPORT_11_en = handshaked & _GEN_1419;
  assign rf_matrix_b_6_tile_v_3_MPORT_11_addr = 8'h53;
  assign rf_matrix_b_6_tile_v_3_MPORT_11_data = rf[rf_matrix_b_6_tile_v_3_MPORT_11_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_6_tile_v_2_MPORT_11_en = handshaked & _GEN_1419;
  assign rf_matrix_b_6_tile_v_2_MPORT_11_addr = 8'h57;
  assign rf_matrix_b_6_tile_v_2_MPORT_11_data = rf[rf_matrix_b_6_tile_v_2_MPORT_11_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_6_tile_v_1_MPORT_11_en = handshaked & _GEN_1419;
  assign rf_matrix_b_6_tile_v_1_MPORT_11_addr = 8'h5b;
  assign rf_matrix_b_6_tile_v_1_MPORT_11_data = rf[rf_matrix_b_6_tile_v_1_MPORT_11_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_6_tile_v_0_MPORT_11_en = handshaked & _GEN_1419;
  assign rf_matrix_b_6_tile_v_0_MPORT_11_addr = 8'h5f;
  assign rf_matrix_b_6_tile_v_0_MPORT_11_data = rf[rf_matrix_b_6_tile_v_0_MPORT_11_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_6_tile_v_3_MPORT_11_en = handshaked & _GEN_1419;
  assign rf_matrix_c_6_tile_v_3_MPORT_11_addr = 8'hb6;
  assign rf_matrix_c_6_tile_v_3_MPORT_11_data = rf[rf_matrix_c_6_tile_v_3_MPORT_11_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_6_tile_v_2_MPORT_11_en = handshaked & _GEN_1419;
  assign rf_matrix_c_6_tile_v_2_MPORT_11_addr = 8'hb7;
  assign rf_matrix_c_6_tile_v_2_MPORT_11_data = rf[rf_matrix_c_6_tile_v_2_MPORT_11_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_6_tile_v_1_MPORT_11_en = handshaked & _GEN_1419;
  assign rf_matrix_c_6_tile_v_1_MPORT_11_addr = 8'hbe;
  assign rf_matrix_c_6_tile_v_1_MPORT_11_data = rf[rf_matrix_c_6_tile_v_1_MPORT_11_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_6_tile_v_0_MPORT_11_en = handshaked & _GEN_1419;
  assign rf_matrix_c_6_tile_v_0_MPORT_11_addr = 8'hbf;
  assign rf_matrix_c_6_tile_v_0_MPORT_11_data = rf[rf_matrix_c_6_tile_v_0_MPORT_11_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_1_MPORT_156_en = handshaked & _GEN_1431;
  assign rf_a_tile_v_1_MPORT_156_addr = 8'h12;
  assign rf_a_tile_v_1_MPORT_156_data = rf[rf_a_tile_v_1_MPORT_156_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_0_MPORT_156_en = handshaked & _GEN_1431;
  assign rf_a_tile_v_0_MPORT_156_addr = 8'h16;
  assign rf_a_tile_v_0_MPORT_156_data = rf[rf_a_tile_v_0_MPORT_156_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_6_tile_v_3_MPORT_12_en = handshaked & _GEN_1431;
  assign rf_matrix_b_6_tile_v_3_MPORT_12_addr = 8'h63;
  assign rf_matrix_b_6_tile_v_3_MPORT_12_data = rf[rf_matrix_b_6_tile_v_3_MPORT_12_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_6_tile_v_2_MPORT_12_en = handshaked & _GEN_1431;
  assign rf_matrix_b_6_tile_v_2_MPORT_12_addr = 8'h67;
  assign rf_matrix_b_6_tile_v_2_MPORT_12_data = rf[rf_matrix_b_6_tile_v_2_MPORT_12_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_6_tile_v_1_MPORT_12_en = handshaked & _GEN_1431;
  assign rf_matrix_b_6_tile_v_1_MPORT_12_addr = 8'h6b;
  assign rf_matrix_b_6_tile_v_1_MPORT_12_data = rf[rf_matrix_b_6_tile_v_1_MPORT_12_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_6_tile_v_0_MPORT_12_en = handshaked & _GEN_1431;
  assign rf_matrix_b_6_tile_v_0_MPORT_12_addr = 8'h6f;
  assign rf_matrix_b_6_tile_v_0_MPORT_12_data = rf[rf_matrix_b_6_tile_v_0_MPORT_12_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_6_tile_v_3_MPORT_12_en = handshaked & _GEN_1431;
  assign rf_matrix_c_6_tile_v_3_MPORT_12_addr = 8'ha4;
  assign rf_matrix_c_6_tile_v_3_MPORT_12_data = rf[rf_matrix_c_6_tile_v_3_MPORT_12_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_6_tile_v_2_MPORT_12_en = handshaked & _GEN_1431;
  assign rf_matrix_c_6_tile_v_2_MPORT_12_addr = 8'ha5;
  assign rf_matrix_c_6_tile_v_2_MPORT_12_data = rf[rf_matrix_c_6_tile_v_2_MPORT_12_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_6_tile_v_1_MPORT_12_en = handshaked & _GEN_1431;
  assign rf_matrix_c_6_tile_v_1_MPORT_12_addr = 8'hac;
  assign rf_matrix_c_6_tile_v_1_MPORT_12_data = rf[rf_matrix_c_6_tile_v_1_MPORT_12_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_6_tile_v_0_MPORT_12_en = handshaked & _GEN_1431;
  assign rf_matrix_c_6_tile_v_0_MPORT_12_addr = 8'had;
  assign rf_matrix_c_6_tile_v_0_MPORT_12_data = rf[rf_matrix_c_6_tile_v_0_MPORT_12_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_3_MPORT_52_en = handshaked & _GEN_1443;
  assign rf_a_tile_v_3_MPORT_52_addr = 8'h12;
  assign rf_a_tile_v_3_MPORT_52_data = rf[rf_a_tile_v_3_MPORT_52_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_2_MPORT_52_en = handshaked & _GEN_1443;
  assign rf_a_tile_v_2_MPORT_52_addr = 8'h16;
  assign rf_a_tile_v_2_MPORT_52_data = rf[rf_a_tile_v_2_MPORT_52_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_1_MPORT_157_en = handshaked & _GEN_1443;
  assign rf_a_tile_v_1_MPORT_157_addr = 8'h1a;
  assign rf_a_tile_v_1_MPORT_157_data = rf[rf_a_tile_v_1_MPORT_157_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_0_MPORT_157_en = handshaked & _GEN_1443;
  assign rf_a_tile_v_0_MPORT_157_addr = 8'h1e;
  assign rf_a_tile_v_0_MPORT_157_data = rf[rf_a_tile_v_0_MPORT_157_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_6_tile_v_3_MPORT_13_en = handshaked & _GEN_1443;
  assign rf_matrix_b_6_tile_v_3_MPORT_13_addr = 8'h63;
  assign rf_matrix_b_6_tile_v_3_MPORT_13_data = rf[rf_matrix_b_6_tile_v_3_MPORT_13_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_6_tile_v_2_MPORT_13_en = handshaked & _GEN_1443;
  assign rf_matrix_b_6_tile_v_2_MPORT_13_addr = 8'h67;
  assign rf_matrix_b_6_tile_v_2_MPORT_13_data = rf[rf_matrix_b_6_tile_v_2_MPORT_13_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_6_tile_v_1_MPORT_13_en = handshaked & _GEN_1443;
  assign rf_matrix_b_6_tile_v_1_MPORT_13_addr = 8'h6b;
  assign rf_matrix_b_6_tile_v_1_MPORT_13_data = rf[rf_matrix_b_6_tile_v_1_MPORT_13_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_6_tile_v_0_MPORT_13_en = handshaked & _GEN_1443;
  assign rf_matrix_b_6_tile_v_0_MPORT_13_addr = 8'h6f;
  assign rf_matrix_b_6_tile_v_0_MPORT_13_data = rf[rf_matrix_b_6_tile_v_0_MPORT_13_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_6_tile_v_3_MPORT_13_en = handshaked & _GEN_1443;
  assign rf_matrix_c_6_tile_v_3_MPORT_13_addr = 8'h92;
  assign rf_matrix_c_6_tile_v_3_MPORT_13_data = rf[rf_matrix_c_6_tile_v_3_MPORT_13_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_6_tile_v_2_MPORT_13_en = handshaked & _GEN_1443;
  assign rf_matrix_c_6_tile_v_2_MPORT_13_addr = 8'h96;
  assign rf_matrix_c_6_tile_v_2_MPORT_13_data = rf[rf_matrix_c_6_tile_v_2_MPORT_13_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_6_tile_v_1_MPORT_13_en = handshaked & _GEN_1443;
  assign rf_matrix_c_6_tile_v_1_MPORT_13_addr = 8'h9a;
  assign rf_matrix_c_6_tile_v_1_MPORT_13_data = rf[rf_matrix_c_6_tile_v_1_MPORT_13_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_6_tile_v_0_MPORT_13_en = handshaked & _GEN_1443;
  assign rf_matrix_c_6_tile_v_0_MPORT_13_addr = 8'h9e;
  assign rf_matrix_c_6_tile_v_0_MPORT_13_data = rf[rf_matrix_c_6_tile_v_0_MPORT_13_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_1_MPORT_158_en = handshaked & _GEN_1457;
  assign rf_a_tile_v_1_MPORT_158_addr = 8'h1a;
  assign rf_a_tile_v_1_MPORT_158_data = rf[rf_a_tile_v_1_MPORT_158_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_0_MPORT_158_en = handshaked & _GEN_1457;
  assign rf_a_tile_v_0_MPORT_158_addr = 8'h1e;
  assign rf_a_tile_v_0_MPORT_158_data = rf[rf_a_tile_v_0_MPORT_158_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_6_tile_v_3_MPORT_14_en = handshaked & _GEN_1457;
  assign rf_matrix_b_6_tile_v_3_MPORT_14_addr = 8'h63;
  assign rf_matrix_b_6_tile_v_3_MPORT_14_data = rf[rf_matrix_b_6_tile_v_3_MPORT_14_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_6_tile_v_2_MPORT_14_en = handshaked & _GEN_1457;
  assign rf_matrix_b_6_tile_v_2_MPORT_14_addr = 8'h67;
  assign rf_matrix_b_6_tile_v_2_MPORT_14_data = rf[rf_matrix_b_6_tile_v_2_MPORT_14_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_6_tile_v_1_MPORT_14_en = handshaked & _GEN_1457;
  assign rf_matrix_b_6_tile_v_1_MPORT_14_addr = 8'h6b;
  assign rf_matrix_b_6_tile_v_1_MPORT_14_data = rf[rf_matrix_b_6_tile_v_1_MPORT_14_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_6_tile_v_0_MPORT_14_en = handshaked & _GEN_1457;
  assign rf_matrix_b_6_tile_v_0_MPORT_14_addr = 8'h6f;
  assign rf_matrix_b_6_tile_v_0_MPORT_14_data = rf[rf_matrix_b_6_tile_v_0_MPORT_14_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_6_tile_v_3_MPORT_14_en = handshaked & _GEN_1457;
  assign rf_matrix_c_6_tile_v_3_MPORT_14_addr = 8'hb4;
  assign rf_matrix_c_6_tile_v_3_MPORT_14_data = rf[rf_matrix_c_6_tile_v_3_MPORT_14_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_6_tile_v_2_MPORT_14_en = handshaked & _GEN_1457;
  assign rf_matrix_c_6_tile_v_2_MPORT_14_addr = 8'hb5;
  assign rf_matrix_c_6_tile_v_2_MPORT_14_data = rf[rf_matrix_c_6_tile_v_2_MPORT_14_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_6_tile_v_1_MPORT_14_en = handshaked & _GEN_1457;
  assign rf_matrix_c_6_tile_v_1_MPORT_14_addr = 8'hbc;
  assign rf_matrix_c_6_tile_v_1_MPORT_14_data = rf[rf_matrix_c_6_tile_v_1_MPORT_14_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_6_tile_v_0_MPORT_14_en = handshaked & _GEN_1457;
  assign rf_matrix_c_6_tile_v_0_MPORT_14_addr = 8'hbd;
  assign rf_matrix_c_6_tile_v_0_MPORT_14_data = rf[rf_matrix_c_6_tile_v_0_MPORT_14_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_3_MPORT_53_en = handshaked & _GEN_1469;
  assign rf_a_tile_v_3_MPORT_53_addr = 8'h12;
  assign rf_a_tile_v_3_MPORT_53_data = rf[rf_a_tile_v_3_MPORT_53_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_2_MPORT_53_en = handshaked & _GEN_1469;
  assign rf_a_tile_v_2_MPORT_53_addr = 8'h16;
  assign rf_a_tile_v_2_MPORT_53_data = rf[rf_a_tile_v_2_MPORT_53_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_1_MPORT_159_en = handshaked & _GEN_1469;
  assign rf_a_tile_v_1_MPORT_159_addr = 8'h1a;
  assign rf_a_tile_v_1_MPORT_159_data = rf[rf_a_tile_v_1_MPORT_159_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_0_MPORT_159_en = handshaked & _GEN_1469;
  assign rf_a_tile_v_0_MPORT_159_addr = 8'h1e;
  assign rf_a_tile_v_0_MPORT_159_data = rf[rf_a_tile_v_0_MPORT_159_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_6_tile_v_3_MPORT_15_en = handshaked & _GEN_1469;
  assign rf_matrix_b_6_tile_v_3_MPORT_15_addr = 8'h63;
  assign rf_matrix_b_6_tile_v_3_MPORT_15_data = rf[rf_matrix_b_6_tile_v_3_MPORT_15_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_6_tile_v_2_MPORT_15_en = handshaked & _GEN_1469;
  assign rf_matrix_b_6_tile_v_2_MPORT_15_addr = 8'h67;
  assign rf_matrix_b_6_tile_v_2_MPORT_15_data = rf[rf_matrix_b_6_tile_v_2_MPORT_15_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_6_tile_v_1_MPORT_15_en = handshaked & _GEN_1469;
  assign rf_matrix_b_6_tile_v_1_MPORT_15_addr = 8'h6b;
  assign rf_matrix_b_6_tile_v_1_MPORT_15_data = rf[rf_matrix_b_6_tile_v_1_MPORT_15_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_6_tile_v_0_MPORT_15_en = handshaked & _GEN_1469;
  assign rf_matrix_b_6_tile_v_0_MPORT_15_addr = 8'h6f;
  assign rf_matrix_b_6_tile_v_0_MPORT_15_data = rf[rf_matrix_b_6_tile_v_0_MPORT_15_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_6_tile_v_3_MPORT_15_en = handshaked & _GEN_1469;
  assign rf_matrix_c_6_tile_v_3_MPORT_15_addr = 8'h93;
  assign rf_matrix_c_6_tile_v_3_MPORT_15_data = rf[rf_matrix_c_6_tile_v_3_MPORT_15_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_6_tile_v_2_MPORT_15_en = handshaked & _GEN_1469;
  assign rf_matrix_c_6_tile_v_2_MPORT_15_addr = 8'h97;
  assign rf_matrix_c_6_tile_v_2_MPORT_15_data = rf[rf_matrix_c_6_tile_v_2_MPORT_15_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_6_tile_v_1_MPORT_15_en = handshaked & _GEN_1469;
  assign rf_matrix_c_6_tile_v_1_MPORT_15_addr = 8'h9b;
  assign rf_matrix_c_6_tile_v_1_MPORT_15_data = rf[rf_matrix_c_6_tile_v_1_MPORT_15_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_6_tile_v_0_MPORT_15_en = handshaked & _GEN_1469;
  assign rf_matrix_c_6_tile_v_0_MPORT_15_addr = 8'h9f;
  assign rf_matrix_c_6_tile_v_0_MPORT_15_data = rf[rf_matrix_c_6_tile_v_0_MPORT_15_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_1_MPORT_160_en = handshaked & _GEN_1483;
  assign rf_a_tile_v_1_MPORT_160_addr = 8'h12;
  assign rf_a_tile_v_1_MPORT_160_data = rf[rf_a_tile_v_1_MPORT_160_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_0_MPORT_160_en = handshaked & _GEN_1483;
  assign rf_a_tile_v_0_MPORT_160_addr = 8'h16;
  assign rf_a_tile_v_0_MPORT_160_data = rf[rf_a_tile_v_0_MPORT_160_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_6_tile_v_3_MPORT_16_en = handshaked & _GEN_1483;
  assign rf_matrix_b_6_tile_v_3_MPORT_16_addr = 8'h63;
  assign rf_matrix_b_6_tile_v_3_MPORT_16_data = rf[rf_matrix_b_6_tile_v_3_MPORT_16_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_6_tile_v_2_MPORT_16_en = handshaked & _GEN_1483;
  assign rf_matrix_b_6_tile_v_2_MPORT_16_addr = 8'h67;
  assign rf_matrix_b_6_tile_v_2_MPORT_16_data = rf[rf_matrix_b_6_tile_v_2_MPORT_16_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_6_tile_v_1_MPORT_16_en = handshaked & _GEN_1483;
  assign rf_matrix_b_6_tile_v_1_MPORT_16_addr = 8'h6b;
  assign rf_matrix_b_6_tile_v_1_MPORT_16_data = rf[rf_matrix_b_6_tile_v_1_MPORT_16_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_6_tile_v_0_MPORT_16_en = handshaked & _GEN_1483;
  assign rf_matrix_b_6_tile_v_0_MPORT_16_addr = 8'h6f;
  assign rf_matrix_b_6_tile_v_0_MPORT_16_data = rf[rf_matrix_b_6_tile_v_0_MPORT_16_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_6_tile_v_3_MPORT_16_en = handshaked & _GEN_1483;
  assign rf_matrix_c_6_tile_v_3_MPORT_16_addr = 8'ha6;
  assign rf_matrix_c_6_tile_v_3_MPORT_16_data = rf[rf_matrix_c_6_tile_v_3_MPORT_16_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_6_tile_v_2_MPORT_16_en = handshaked & _GEN_1483;
  assign rf_matrix_c_6_tile_v_2_MPORT_16_addr = 8'ha7;
  assign rf_matrix_c_6_tile_v_2_MPORT_16_data = rf[rf_matrix_c_6_tile_v_2_MPORT_16_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_6_tile_v_1_MPORT_16_en = handshaked & _GEN_1483;
  assign rf_matrix_c_6_tile_v_1_MPORT_16_addr = 8'hae;
  assign rf_matrix_c_6_tile_v_1_MPORT_16_data = rf[rf_matrix_c_6_tile_v_1_MPORT_16_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_6_tile_v_0_MPORT_16_en = handshaked & _GEN_1483;
  assign rf_matrix_c_6_tile_v_0_MPORT_16_addr = 8'haf;
  assign rf_matrix_c_6_tile_v_0_MPORT_16_data = rf[rf_matrix_c_6_tile_v_0_MPORT_16_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_1_MPORT_161_en = handshaked & _GEN_1495;
  assign rf_a_tile_v_1_MPORT_161_addr = 8'h1a;
  assign rf_a_tile_v_1_MPORT_161_data = rf[rf_a_tile_v_1_MPORT_161_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_0_MPORT_161_en = handshaked & _GEN_1495;
  assign rf_a_tile_v_0_MPORT_161_addr = 8'h1e;
  assign rf_a_tile_v_0_MPORT_161_data = rf[rf_a_tile_v_0_MPORT_161_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_6_tile_v_3_MPORT_17_en = handshaked & _GEN_1495;
  assign rf_matrix_b_6_tile_v_3_MPORT_17_addr = 8'h63;
  assign rf_matrix_b_6_tile_v_3_MPORT_17_data = rf[rf_matrix_b_6_tile_v_3_MPORT_17_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_6_tile_v_2_MPORT_17_en = handshaked & _GEN_1495;
  assign rf_matrix_b_6_tile_v_2_MPORT_17_addr = 8'h67;
  assign rf_matrix_b_6_tile_v_2_MPORT_17_data = rf[rf_matrix_b_6_tile_v_2_MPORT_17_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_6_tile_v_1_MPORT_17_en = handshaked & _GEN_1495;
  assign rf_matrix_b_6_tile_v_1_MPORT_17_addr = 8'h6b;
  assign rf_matrix_b_6_tile_v_1_MPORT_17_data = rf[rf_matrix_b_6_tile_v_1_MPORT_17_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_6_tile_v_0_MPORT_17_en = handshaked & _GEN_1495;
  assign rf_matrix_b_6_tile_v_0_MPORT_17_addr = 8'h6f;
  assign rf_matrix_b_6_tile_v_0_MPORT_17_data = rf[rf_matrix_b_6_tile_v_0_MPORT_17_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_6_tile_v_3_MPORT_17_en = handshaked & _GEN_1495;
  assign rf_matrix_c_6_tile_v_3_MPORT_17_addr = 8'hb6;
  assign rf_matrix_c_6_tile_v_3_MPORT_17_data = rf[rf_matrix_c_6_tile_v_3_MPORT_17_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_6_tile_v_2_MPORT_17_en = handshaked & _GEN_1495;
  assign rf_matrix_c_6_tile_v_2_MPORT_17_addr = 8'hb7;
  assign rf_matrix_c_6_tile_v_2_MPORT_17_data = rf[rf_matrix_c_6_tile_v_2_MPORT_17_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_6_tile_v_1_MPORT_17_en = handshaked & _GEN_1495;
  assign rf_matrix_c_6_tile_v_1_MPORT_17_addr = 8'hbe;
  assign rf_matrix_c_6_tile_v_1_MPORT_17_data = rf[rf_matrix_c_6_tile_v_1_MPORT_17_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_6_tile_v_0_MPORT_17_en = handshaked & _GEN_1495;
  assign rf_matrix_c_6_tile_v_0_MPORT_17_addr = 8'hbf;
  assign rf_matrix_c_6_tile_v_0_MPORT_17_data = rf[rf_matrix_c_6_tile_v_0_MPORT_17_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_1_MPORT_162_en = handshaked & _GEN_1507;
  assign rf_a_tile_v_1_MPORT_162_addr = 8'h13;
  assign rf_a_tile_v_1_MPORT_162_data = rf[rf_a_tile_v_1_MPORT_162_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_0_MPORT_162_en = handshaked & _GEN_1507;
  assign rf_a_tile_v_0_MPORT_162_addr = 8'h17;
  assign rf_a_tile_v_0_MPORT_162_data = rf[rf_a_tile_v_0_MPORT_162_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_6_tile_v_3_MPORT_18_en = handshaked & _GEN_1507;
  assign rf_matrix_b_6_tile_v_3_MPORT_18_addr = 8'h73;
  assign rf_matrix_b_6_tile_v_3_MPORT_18_data = rf[rf_matrix_b_6_tile_v_3_MPORT_18_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_6_tile_v_2_MPORT_18_en = handshaked & _GEN_1507;
  assign rf_matrix_b_6_tile_v_2_MPORT_18_addr = 8'h77;
  assign rf_matrix_b_6_tile_v_2_MPORT_18_data = rf[rf_matrix_b_6_tile_v_2_MPORT_18_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_6_tile_v_1_MPORT_18_en = handshaked & _GEN_1507;
  assign rf_matrix_b_6_tile_v_1_MPORT_18_addr = 8'h7b;
  assign rf_matrix_b_6_tile_v_1_MPORT_18_data = rf[rf_matrix_b_6_tile_v_1_MPORT_18_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_6_tile_v_0_MPORT_18_en = handshaked & _GEN_1507;
  assign rf_matrix_b_6_tile_v_0_MPORT_18_addr = 8'h7f;
  assign rf_matrix_b_6_tile_v_0_MPORT_18_data = rf[rf_matrix_b_6_tile_v_0_MPORT_18_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_6_tile_v_3_MPORT_18_en = handshaked & _GEN_1507;
  assign rf_matrix_c_6_tile_v_3_MPORT_18_addr = 8'ha4;
  assign rf_matrix_c_6_tile_v_3_MPORT_18_data = rf[rf_matrix_c_6_tile_v_3_MPORT_18_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_6_tile_v_2_MPORT_18_en = handshaked & _GEN_1507;
  assign rf_matrix_c_6_tile_v_2_MPORT_18_addr = 8'ha5;
  assign rf_matrix_c_6_tile_v_2_MPORT_18_data = rf[rf_matrix_c_6_tile_v_2_MPORT_18_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_6_tile_v_1_MPORT_18_en = handshaked & _GEN_1507;
  assign rf_matrix_c_6_tile_v_1_MPORT_18_addr = 8'hac;
  assign rf_matrix_c_6_tile_v_1_MPORT_18_data = rf[rf_matrix_c_6_tile_v_1_MPORT_18_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_6_tile_v_0_MPORT_18_en = handshaked & _GEN_1507;
  assign rf_matrix_c_6_tile_v_0_MPORT_18_addr = 8'had;
  assign rf_matrix_c_6_tile_v_0_MPORT_18_data = rf[rf_matrix_c_6_tile_v_0_MPORT_18_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_3_MPORT_54_en = handshaked & _GEN_1519;
  assign rf_a_tile_v_3_MPORT_54_addr = 8'h13;
  assign rf_a_tile_v_3_MPORT_54_data = rf[rf_a_tile_v_3_MPORT_54_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_2_MPORT_54_en = handshaked & _GEN_1519;
  assign rf_a_tile_v_2_MPORT_54_addr = 8'h17;
  assign rf_a_tile_v_2_MPORT_54_data = rf[rf_a_tile_v_2_MPORT_54_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_1_MPORT_163_en = handshaked & _GEN_1519;
  assign rf_a_tile_v_1_MPORT_163_addr = 8'h1b;
  assign rf_a_tile_v_1_MPORT_163_data = rf[rf_a_tile_v_1_MPORT_163_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_0_MPORT_163_en = handshaked & _GEN_1519;
  assign rf_a_tile_v_0_MPORT_163_addr = 8'h1f;
  assign rf_a_tile_v_0_MPORT_163_data = rf[rf_a_tile_v_0_MPORT_163_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_6_tile_v_3_MPORT_19_en = handshaked & _GEN_1519;
  assign rf_matrix_b_6_tile_v_3_MPORT_19_addr = 8'h73;
  assign rf_matrix_b_6_tile_v_3_MPORT_19_data = rf[rf_matrix_b_6_tile_v_3_MPORT_19_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_6_tile_v_2_MPORT_19_en = handshaked & _GEN_1519;
  assign rf_matrix_b_6_tile_v_2_MPORT_19_addr = 8'h77;
  assign rf_matrix_b_6_tile_v_2_MPORT_19_data = rf[rf_matrix_b_6_tile_v_2_MPORT_19_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_6_tile_v_1_MPORT_19_en = handshaked & _GEN_1519;
  assign rf_matrix_b_6_tile_v_1_MPORT_19_addr = 8'h7b;
  assign rf_matrix_b_6_tile_v_1_MPORT_19_data = rf[rf_matrix_b_6_tile_v_1_MPORT_19_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_6_tile_v_0_MPORT_19_en = handshaked & _GEN_1519;
  assign rf_matrix_b_6_tile_v_0_MPORT_19_addr = 8'h7f;
  assign rf_matrix_b_6_tile_v_0_MPORT_19_data = rf[rf_matrix_b_6_tile_v_0_MPORT_19_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_6_tile_v_3_MPORT_19_en = handshaked & _GEN_1519;
  assign rf_matrix_c_6_tile_v_3_MPORT_19_addr = 8'h92;
  assign rf_matrix_c_6_tile_v_3_MPORT_19_data = rf[rf_matrix_c_6_tile_v_3_MPORT_19_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_6_tile_v_2_MPORT_19_en = handshaked & _GEN_1519;
  assign rf_matrix_c_6_tile_v_2_MPORT_19_addr = 8'h96;
  assign rf_matrix_c_6_tile_v_2_MPORT_19_data = rf[rf_matrix_c_6_tile_v_2_MPORT_19_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_6_tile_v_1_MPORT_19_en = handshaked & _GEN_1519;
  assign rf_matrix_c_6_tile_v_1_MPORT_19_addr = 8'h9a;
  assign rf_matrix_c_6_tile_v_1_MPORT_19_data = rf[rf_matrix_c_6_tile_v_1_MPORT_19_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_6_tile_v_0_MPORT_19_en = handshaked & _GEN_1519;
  assign rf_matrix_c_6_tile_v_0_MPORT_19_addr = 8'h9e;
  assign rf_matrix_c_6_tile_v_0_MPORT_19_data = rf[rf_matrix_c_6_tile_v_0_MPORT_19_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_1_MPORT_164_en = handshaked & _GEN_1533;
  assign rf_a_tile_v_1_MPORT_164_addr = 8'h1b;
  assign rf_a_tile_v_1_MPORT_164_data = rf[rf_a_tile_v_1_MPORT_164_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_0_MPORT_164_en = handshaked & _GEN_1533;
  assign rf_a_tile_v_0_MPORT_164_addr = 8'h1f;
  assign rf_a_tile_v_0_MPORT_164_data = rf[rf_a_tile_v_0_MPORT_164_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_6_tile_v_3_MPORT_20_en = handshaked & _GEN_1533;
  assign rf_matrix_b_6_tile_v_3_MPORT_20_addr = 8'h73;
  assign rf_matrix_b_6_tile_v_3_MPORT_20_data = rf[rf_matrix_b_6_tile_v_3_MPORT_20_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_6_tile_v_2_MPORT_20_en = handshaked & _GEN_1533;
  assign rf_matrix_b_6_tile_v_2_MPORT_20_addr = 8'h77;
  assign rf_matrix_b_6_tile_v_2_MPORT_20_data = rf[rf_matrix_b_6_tile_v_2_MPORT_20_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_6_tile_v_1_MPORT_20_en = handshaked & _GEN_1533;
  assign rf_matrix_b_6_tile_v_1_MPORT_20_addr = 8'h7b;
  assign rf_matrix_b_6_tile_v_1_MPORT_20_data = rf[rf_matrix_b_6_tile_v_1_MPORT_20_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_6_tile_v_0_MPORT_20_en = handshaked & _GEN_1533;
  assign rf_matrix_b_6_tile_v_0_MPORT_20_addr = 8'h7f;
  assign rf_matrix_b_6_tile_v_0_MPORT_20_data = rf[rf_matrix_b_6_tile_v_0_MPORT_20_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_6_tile_v_3_MPORT_20_en = handshaked & _GEN_1533;
  assign rf_matrix_c_6_tile_v_3_MPORT_20_addr = 8'hb4;
  assign rf_matrix_c_6_tile_v_3_MPORT_20_data = rf[rf_matrix_c_6_tile_v_3_MPORT_20_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_6_tile_v_2_MPORT_20_en = handshaked & _GEN_1533;
  assign rf_matrix_c_6_tile_v_2_MPORT_20_addr = 8'hb5;
  assign rf_matrix_c_6_tile_v_2_MPORT_20_data = rf[rf_matrix_c_6_tile_v_2_MPORT_20_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_6_tile_v_1_MPORT_20_en = handshaked & _GEN_1533;
  assign rf_matrix_c_6_tile_v_1_MPORT_20_addr = 8'hbc;
  assign rf_matrix_c_6_tile_v_1_MPORT_20_data = rf[rf_matrix_c_6_tile_v_1_MPORT_20_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_6_tile_v_0_MPORT_20_en = handshaked & _GEN_1533;
  assign rf_matrix_c_6_tile_v_0_MPORT_20_addr = 8'hbd;
  assign rf_matrix_c_6_tile_v_0_MPORT_20_data = rf[rf_matrix_c_6_tile_v_0_MPORT_20_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_3_MPORT_55_en = handshaked & _GEN_1545;
  assign rf_a_tile_v_3_MPORT_55_addr = 8'h13;
  assign rf_a_tile_v_3_MPORT_55_data = rf[rf_a_tile_v_3_MPORT_55_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_2_MPORT_55_en = handshaked & _GEN_1545;
  assign rf_a_tile_v_2_MPORT_55_addr = 8'h17;
  assign rf_a_tile_v_2_MPORT_55_data = rf[rf_a_tile_v_2_MPORT_55_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_1_MPORT_165_en = handshaked & _GEN_1545;
  assign rf_a_tile_v_1_MPORT_165_addr = 8'h1b;
  assign rf_a_tile_v_1_MPORT_165_data = rf[rf_a_tile_v_1_MPORT_165_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_0_MPORT_165_en = handshaked & _GEN_1545;
  assign rf_a_tile_v_0_MPORT_165_addr = 8'h1f;
  assign rf_a_tile_v_0_MPORT_165_data = rf[rf_a_tile_v_0_MPORT_165_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_6_tile_v_3_MPORT_21_en = handshaked & _GEN_1545;
  assign rf_matrix_b_6_tile_v_3_MPORT_21_addr = 8'h73;
  assign rf_matrix_b_6_tile_v_3_MPORT_21_data = rf[rf_matrix_b_6_tile_v_3_MPORT_21_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_6_tile_v_2_MPORT_21_en = handshaked & _GEN_1545;
  assign rf_matrix_b_6_tile_v_2_MPORT_21_addr = 8'h77;
  assign rf_matrix_b_6_tile_v_2_MPORT_21_data = rf[rf_matrix_b_6_tile_v_2_MPORT_21_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_6_tile_v_1_MPORT_21_en = handshaked & _GEN_1545;
  assign rf_matrix_b_6_tile_v_1_MPORT_21_addr = 8'h7b;
  assign rf_matrix_b_6_tile_v_1_MPORT_21_data = rf[rf_matrix_b_6_tile_v_1_MPORT_21_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_6_tile_v_0_MPORT_21_en = handshaked & _GEN_1545;
  assign rf_matrix_b_6_tile_v_0_MPORT_21_addr = 8'h7f;
  assign rf_matrix_b_6_tile_v_0_MPORT_21_data = rf[rf_matrix_b_6_tile_v_0_MPORT_21_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_6_tile_v_3_MPORT_21_en = handshaked & _GEN_1545;
  assign rf_matrix_c_6_tile_v_3_MPORT_21_addr = 8'h93;
  assign rf_matrix_c_6_tile_v_3_MPORT_21_data = rf[rf_matrix_c_6_tile_v_3_MPORT_21_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_6_tile_v_2_MPORT_21_en = handshaked & _GEN_1545;
  assign rf_matrix_c_6_tile_v_2_MPORT_21_addr = 8'h97;
  assign rf_matrix_c_6_tile_v_2_MPORT_21_data = rf[rf_matrix_c_6_tile_v_2_MPORT_21_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_6_tile_v_1_MPORT_21_en = handshaked & _GEN_1545;
  assign rf_matrix_c_6_tile_v_1_MPORT_21_addr = 8'h9b;
  assign rf_matrix_c_6_tile_v_1_MPORT_21_data = rf[rf_matrix_c_6_tile_v_1_MPORT_21_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_6_tile_v_0_MPORT_21_en = handshaked & _GEN_1545;
  assign rf_matrix_c_6_tile_v_0_MPORT_21_addr = 8'h9f;
  assign rf_matrix_c_6_tile_v_0_MPORT_21_data = rf[rf_matrix_c_6_tile_v_0_MPORT_21_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_1_MPORT_166_en = handshaked & _GEN_1559;
  assign rf_a_tile_v_1_MPORT_166_addr = 8'h13;
  assign rf_a_tile_v_1_MPORT_166_data = rf[rf_a_tile_v_1_MPORT_166_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_0_MPORT_166_en = handshaked & _GEN_1559;
  assign rf_a_tile_v_0_MPORT_166_addr = 8'h17;
  assign rf_a_tile_v_0_MPORT_166_data = rf[rf_a_tile_v_0_MPORT_166_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_6_tile_v_3_MPORT_22_en = handshaked & _GEN_1559;
  assign rf_matrix_b_6_tile_v_3_MPORT_22_addr = 8'h73;
  assign rf_matrix_b_6_tile_v_3_MPORT_22_data = rf[rf_matrix_b_6_tile_v_3_MPORT_22_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_6_tile_v_2_MPORT_22_en = handshaked & _GEN_1559;
  assign rf_matrix_b_6_tile_v_2_MPORT_22_addr = 8'h77;
  assign rf_matrix_b_6_tile_v_2_MPORT_22_data = rf[rf_matrix_b_6_tile_v_2_MPORT_22_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_6_tile_v_1_MPORT_22_en = handshaked & _GEN_1559;
  assign rf_matrix_b_6_tile_v_1_MPORT_22_addr = 8'h7b;
  assign rf_matrix_b_6_tile_v_1_MPORT_22_data = rf[rf_matrix_b_6_tile_v_1_MPORT_22_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_6_tile_v_0_MPORT_22_en = handshaked & _GEN_1559;
  assign rf_matrix_b_6_tile_v_0_MPORT_22_addr = 8'h7f;
  assign rf_matrix_b_6_tile_v_0_MPORT_22_data = rf[rf_matrix_b_6_tile_v_0_MPORT_22_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_6_tile_v_3_MPORT_22_en = handshaked & _GEN_1559;
  assign rf_matrix_c_6_tile_v_3_MPORT_22_addr = 8'ha6;
  assign rf_matrix_c_6_tile_v_3_MPORT_22_data = rf[rf_matrix_c_6_tile_v_3_MPORT_22_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_6_tile_v_2_MPORT_22_en = handshaked & _GEN_1559;
  assign rf_matrix_c_6_tile_v_2_MPORT_22_addr = 8'ha7;
  assign rf_matrix_c_6_tile_v_2_MPORT_22_data = rf[rf_matrix_c_6_tile_v_2_MPORT_22_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_6_tile_v_1_MPORT_22_en = handshaked & _GEN_1559;
  assign rf_matrix_c_6_tile_v_1_MPORT_22_addr = 8'hae;
  assign rf_matrix_c_6_tile_v_1_MPORT_22_data = rf[rf_matrix_c_6_tile_v_1_MPORT_22_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_6_tile_v_0_MPORT_22_en = handshaked & _GEN_1559;
  assign rf_matrix_c_6_tile_v_0_MPORT_22_addr = 8'haf;
  assign rf_matrix_c_6_tile_v_0_MPORT_22_data = rf[rf_matrix_c_6_tile_v_0_MPORT_22_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_1_MPORT_167_en = handshaked & _GEN_1571;
  assign rf_a_tile_v_1_MPORT_167_addr = 8'h1b;
  assign rf_a_tile_v_1_MPORT_167_data = rf[rf_a_tile_v_1_MPORT_167_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_0_MPORT_167_en = handshaked & _GEN_1571;
  assign rf_a_tile_v_0_MPORT_167_addr = 8'h1f;
  assign rf_a_tile_v_0_MPORT_167_data = rf[rf_a_tile_v_0_MPORT_167_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_6_tile_v_3_MPORT_23_en = handshaked & _GEN_1571;
  assign rf_matrix_b_6_tile_v_3_MPORT_23_addr = 8'h73;
  assign rf_matrix_b_6_tile_v_3_MPORT_23_data = rf[rf_matrix_b_6_tile_v_3_MPORT_23_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_6_tile_v_2_MPORT_23_en = handshaked & _GEN_1571;
  assign rf_matrix_b_6_tile_v_2_MPORT_23_addr = 8'h77;
  assign rf_matrix_b_6_tile_v_2_MPORT_23_data = rf[rf_matrix_b_6_tile_v_2_MPORT_23_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_6_tile_v_1_MPORT_23_en = handshaked & _GEN_1571;
  assign rf_matrix_b_6_tile_v_1_MPORT_23_addr = 8'h7b;
  assign rf_matrix_b_6_tile_v_1_MPORT_23_data = rf[rf_matrix_b_6_tile_v_1_MPORT_23_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_6_tile_v_0_MPORT_23_en = handshaked & _GEN_1571;
  assign rf_matrix_b_6_tile_v_0_MPORT_23_addr = 8'h7f;
  assign rf_matrix_b_6_tile_v_0_MPORT_23_data = rf[rf_matrix_b_6_tile_v_0_MPORT_23_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_6_tile_v_3_MPORT_23_en = handshaked & _GEN_1571;
  assign rf_matrix_c_6_tile_v_3_MPORT_23_addr = 8'hb6;
  assign rf_matrix_c_6_tile_v_3_MPORT_23_data = rf[rf_matrix_c_6_tile_v_3_MPORT_23_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_6_tile_v_2_MPORT_23_en = handshaked & _GEN_1571;
  assign rf_matrix_c_6_tile_v_2_MPORT_23_addr = 8'hb7;
  assign rf_matrix_c_6_tile_v_2_MPORT_23_data = rf[rf_matrix_c_6_tile_v_2_MPORT_23_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_6_tile_v_1_MPORT_23_en = handshaked & _GEN_1571;
  assign rf_matrix_c_6_tile_v_1_MPORT_23_addr = 8'hbe;
  assign rf_matrix_c_6_tile_v_1_MPORT_23_data = rf[rf_matrix_c_6_tile_v_1_MPORT_23_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_6_tile_v_0_MPORT_23_en = handshaked & _GEN_1571;
  assign rf_matrix_c_6_tile_v_0_MPORT_23_addr = 8'hbf;
  assign rf_matrix_c_6_tile_v_0_MPORT_23_data = rf[rf_matrix_c_6_tile_v_0_MPORT_23_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_1_MPORT_168_en = handshaked & _GEN_1276;
  assign rf_a_tile_v_1_MPORT_168_addr = 8'h30;
  assign rf_a_tile_v_1_MPORT_168_data = rf[rf_a_tile_v_1_MPORT_168_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_0_MPORT_168_en = handshaked & _GEN_1276;
  assign rf_a_tile_v_0_MPORT_168_addr = 8'h34;
  assign rf_a_tile_v_0_MPORT_168_data = rf[rf_a_tile_v_0_MPORT_168_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_7_tile_v_3_MPORT_en = handshaked & _GEN_1276;
  assign rf_matrix_b_7_tile_v_3_MPORT_addr = 8'h43;
  assign rf_matrix_b_7_tile_v_3_MPORT_data = rf[rf_matrix_b_7_tile_v_3_MPORT_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_7_tile_v_2_MPORT_en = handshaked & _GEN_1276;
  assign rf_matrix_b_7_tile_v_2_MPORT_addr = 8'h47;
  assign rf_matrix_b_7_tile_v_2_MPORT_data = rf[rf_matrix_b_7_tile_v_2_MPORT_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_7_tile_v_1_MPORT_en = handshaked & _GEN_1276;
  assign rf_matrix_b_7_tile_v_1_MPORT_addr = 8'h4b;
  assign rf_matrix_b_7_tile_v_1_MPORT_data = rf[rf_matrix_b_7_tile_v_1_MPORT_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_7_tile_v_0_MPORT_en = handshaked & _GEN_1276;
  assign rf_matrix_b_7_tile_v_0_MPORT_addr = 8'h4f;
  assign rf_matrix_b_7_tile_v_0_MPORT_data = rf[rf_matrix_b_7_tile_v_0_MPORT_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_7_tile_v_3_MPORT_en = handshaked & _GEN_1276;
  assign rf_matrix_c_7_tile_v_3_MPORT_addr = 8'he4;
  assign rf_matrix_c_7_tile_v_3_MPORT_data = rf[rf_matrix_c_7_tile_v_3_MPORT_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_7_tile_v_2_MPORT_en = handshaked & _GEN_1276;
  assign rf_matrix_c_7_tile_v_2_MPORT_addr = 8'he5;
  assign rf_matrix_c_7_tile_v_2_MPORT_data = rf[rf_matrix_c_7_tile_v_2_MPORT_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_7_tile_v_1_MPORT_en = handshaked & _GEN_1276;
  assign rf_matrix_c_7_tile_v_1_MPORT_addr = 8'hec;
  assign rf_matrix_c_7_tile_v_1_MPORT_data = rf[rf_matrix_c_7_tile_v_1_MPORT_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_7_tile_v_0_MPORT_en = handshaked & _GEN_1276;
  assign rf_matrix_c_7_tile_v_0_MPORT_addr = 8'hed;
  assign rf_matrix_c_7_tile_v_0_MPORT_data = rf[rf_matrix_c_7_tile_v_0_MPORT_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_3_MPORT_56_en = handshaked & _GEN_1291;
  assign rf_a_tile_v_3_MPORT_56_addr = 8'h30;
  assign rf_a_tile_v_3_MPORT_56_data = rf[rf_a_tile_v_3_MPORT_56_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_2_MPORT_56_en = handshaked & _GEN_1291;
  assign rf_a_tile_v_2_MPORT_56_addr = 8'h34;
  assign rf_a_tile_v_2_MPORT_56_data = rf[rf_a_tile_v_2_MPORT_56_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_1_MPORT_169_en = handshaked & _GEN_1291;
  assign rf_a_tile_v_1_MPORT_169_addr = 8'h38;
  assign rf_a_tile_v_1_MPORT_169_data = rf[rf_a_tile_v_1_MPORT_169_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_0_MPORT_169_en = handshaked & _GEN_1291;
  assign rf_a_tile_v_0_MPORT_169_addr = 8'h3c;
  assign rf_a_tile_v_0_MPORT_169_data = rf[rf_a_tile_v_0_MPORT_169_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_7_tile_v_3_MPORT_1_en = handshaked & _GEN_1291;
  assign rf_matrix_b_7_tile_v_3_MPORT_1_addr = 8'h43;
  assign rf_matrix_b_7_tile_v_3_MPORT_1_data = rf[rf_matrix_b_7_tile_v_3_MPORT_1_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_7_tile_v_2_MPORT_1_en = handshaked & _GEN_1291;
  assign rf_matrix_b_7_tile_v_2_MPORT_1_addr = 8'h47;
  assign rf_matrix_b_7_tile_v_2_MPORT_1_data = rf[rf_matrix_b_7_tile_v_2_MPORT_1_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_7_tile_v_1_MPORT_1_en = handshaked & _GEN_1291;
  assign rf_matrix_b_7_tile_v_1_MPORT_1_addr = 8'h4b;
  assign rf_matrix_b_7_tile_v_1_MPORT_1_data = rf[rf_matrix_b_7_tile_v_1_MPORT_1_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_7_tile_v_0_MPORT_1_en = handshaked & _GEN_1291;
  assign rf_matrix_b_7_tile_v_0_MPORT_1_addr = 8'h4f;
  assign rf_matrix_b_7_tile_v_0_MPORT_1_data = rf[rf_matrix_b_7_tile_v_0_MPORT_1_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_7_tile_v_3_MPORT_1_en = handshaked & _GEN_1291;
  assign rf_matrix_c_7_tile_v_3_MPORT_1_addr = 8'hb2;
  assign rf_matrix_c_7_tile_v_3_MPORT_1_data = rf[rf_matrix_c_7_tile_v_3_MPORT_1_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_7_tile_v_2_MPORT_1_en = handshaked & _GEN_1291;
  assign rf_matrix_c_7_tile_v_2_MPORT_1_addr = 8'hb6;
  assign rf_matrix_c_7_tile_v_2_MPORT_1_data = rf[rf_matrix_c_7_tile_v_2_MPORT_1_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_7_tile_v_1_MPORT_1_en = handshaked & _GEN_1291;
  assign rf_matrix_c_7_tile_v_1_MPORT_1_addr = 8'hba;
  assign rf_matrix_c_7_tile_v_1_MPORT_1_data = rf[rf_matrix_c_7_tile_v_1_MPORT_1_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_7_tile_v_0_MPORT_1_en = handshaked & _GEN_1291;
  assign rf_matrix_c_7_tile_v_0_MPORT_1_addr = 8'hbe;
  assign rf_matrix_c_7_tile_v_0_MPORT_1_data = rf[rf_matrix_c_7_tile_v_0_MPORT_1_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_1_MPORT_170_en = handshaked & _GEN_1305;
  assign rf_a_tile_v_1_MPORT_170_addr = 8'h38;
  assign rf_a_tile_v_1_MPORT_170_data = rf[rf_a_tile_v_1_MPORT_170_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_0_MPORT_170_en = handshaked & _GEN_1305;
  assign rf_a_tile_v_0_MPORT_170_addr = 8'h3c;
  assign rf_a_tile_v_0_MPORT_170_data = rf[rf_a_tile_v_0_MPORT_170_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_7_tile_v_3_MPORT_2_en = handshaked & _GEN_1305;
  assign rf_matrix_b_7_tile_v_3_MPORT_2_addr = 8'h43;
  assign rf_matrix_b_7_tile_v_3_MPORT_2_data = rf[rf_matrix_b_7_tile_v_3_MPORT_2_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_7_tile_v_2_MPORT_2_en = handshaked & _GEN_1305;
  assign rf_matrix_b_7_tile_v_2_MPORT_2_addr = 8'h47;
  assign rf_matrix_b_7_tile_v_2_MPORT_2_data = rf[rf_matrix_b_7_tile_v_2_MPORT_2_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_7_tile_v_1_MPORT_2_en = handshaked & _GEN_1305;
  assign rf_matrix_b_7_tile_v_1_MPORT_2_addr = 8'h4b;
  assign rf_matrix_b_7_tile_v_1_MPORT_2_data = rf[rf_matrix_b_7_tile_v_1_MPORT_2_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_7_tile_v_0_MPORT_2_en = handshaked & _GEN_1305;
  assign rf_matrix_b_7_tile_v_0_MPORT_2_addr = 8'h4f;
  assign rf_matrix_b_7_tile_v_0_MPORT_2_data = rf[rf_matrix_b_7_tile_v_0_MPORT_2_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_7_tile_v_3_MPORT_2_en = handshaked & _GEN_1305;
  assign rf_matrix_c_7_tile_v_3_MPORT_2_addr = 8'hf4;
  assign rf_matrix_c_7_tile_v_3_MPORT_2_data = rf[rf_matrix_c_7_tile_v_3_MPORT_2_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_7_tile_v_2_MPORT_2_en = handshaked & _GEN_1305;
  assign rf_matrix_c_7_tile_v_2_MPORT_2_addr = 8'hf5;
  assign rf_matrix_c_7_tile_v_2_MPORT_2_data = rf[rf_matrix_c_7_tile_v_2_MPORT_2_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_7_tile_v_1_MPORT_2_en = handshaked & _GEN_1305;
  assign rf_matrix_c_7_tile_v_1_MPORT_2_addr = 8'hfc;
  assign rf_matrix_c_7_tile_v_1_MPORT_2_data = rf[rf_matrix_c_7_tile_v_1_MPORT_2_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_7_tile_v_0_MPORT_2_en = handshaked & _GEN_1305;
  assign rf_matrix_c_7_tile_v_0_MPORT_2_addr = 8'hfd;
  assign rf_matrix_c_7_tile_v_0_MPORT_2_data = rf[rf_matrix_c_7_tile_v_0_MPORT_2_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_3_MPORT_57_en = handshaked & _GEN_1317;
  assign rf_a_tile_v_3_MPORT_57_addr = 8'h30;
  assign rf_a_tile_v_3_MPORT_57_data = rf[rf_a_tile_v_3_MPORT_57_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_2_MPORT_57_en = handshaked & _GEN_1317;
  assign rf_a_tile_v_2_MPORT_57_addr = 8'h34;
  assign rf_a_tile_v_2_MPORT_57_data = rf[rf_a_tile_v_2_MPORT_57_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_1_MPORT_171_en = handshaked & _GEN_1317;
  assign rf_a_tile_v_1_MPORT_171_addr = 8'h38;
  assign rf_a_tile_v_1_MPORT_171_data = rf[rf_a_tile_v_1_MPORT_171_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_0_MPORT_171_en = handshaked & _GEN_1317;
  assign rf_a_tile_v_0_MPORT_171_addr = 8'h3c;
  assign rf_a_tile_v_0_MPORT_171_data = rf[rf_a_tile_v_0_MPORT_171_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_7_tile_v_3_MPORT_3_en = handshaked & _GEN_1317;
  assign rf_matrix_b_7_tile_v_3_MPORT_3_addr = 8'h43;
  assign rf_matrix_b_7_tile_v_3_MPORT_3_data = rf[rf_matrix_b_7_tile_v_3_MPORT_3_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_7_tile_v_2_MPORT_3_en = handshaked & _GEN_1317;
  assign rf_matrix_b_7_tile_v_2_MPORT_3_addr = 8'h47;
  assign rf_matrix_b_7_tile_v_2_MPORT_3_data = rf[rf_matrix_b_7_tile_v_2_MPORT_3_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_7_tile_v_1_MPORT_3_en = handshaked & _GEN_1317;
  assign rf_matrix_b_7_tile_v_1_MPORT_3_addr = 8'h4b;
  assign rf_matrix_b_7_tile_v_1_MPORT_3_data = rf[rf_matrix_b_7_tile_v_1_MPORT_3_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_7_tile_v_0_MPORT_3_en = handshaked & _GEN_1317;
  assign rf_matrix_b_7_tile_v_0_MPORT_3_addr = 8'h4f;
  assign rf_matrix_b_7_tile_v_0_MPORT_3_data = rf[rf_matrix_b_7_tile_v_0_MPORT_3_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_7_tile_v_3_MPORT_3_en = handshaked & _GEN_1317;
  assign rf_matrix_c_7_tile_v_3_MPORT_3_addr = 8'hb3;
  assign rf_matrix_c_7_tile_v_3_MPORT_3_data = rf[rf_matrix_c_7_tile_v_3_MPORT_3_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_7_tile_v_2_MPORT_3_en = handshaked & _GEN_1317;
  assign rf_matrix_c_7_tile_v_2_MPORT_3_addr = 8'hb7;
  assign rf_matrix_c_7_tile_v_2_MPORT_3_data = rf[rf_matrix_c_7_tile_v_2_MPORT_3_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_7_tile_v_1_MPORT_3_en = handshaked & _GEN_1317;
  assign rf_matrix_c_7_tile_v_1_MPORT_3_addr = 8'hbb;
  assign rf_matrix_c_7_tile_v_1_MPORT_3_data = rf[rf_matrix_c_7_tile_v_1_MPORT_3_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_7_tile_v_0_MPORT_3_en = handshaked & _GEN_1317;
  assign rf_matrix_c_7_tile_v_0_MPORT_3_addr = 8'hbf;
  assign rf_matrix_c_7_tile_v_0_MPORT_3_data = rf[rf_matrix_c_7_tile_v_0_MPORT_3_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_1_MPORT_172_en = handshaked & _GEN_1331;
  assign rf_a_tile_v_1_MPORT_172_addr = 8'h30;
  assign rf_a_tile_v_1_MPORT_172_data = rf[rf_a_tile_v_1_MPORT_172_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_0_MPORT_172_en = handshaked & _GEN_1331;
  assign rf_a_tile_v_0_MPORT_172_addr = 8'h34;
  assign rf_a_tile_v_0_MPORT_172_data = rf[rf_a_tile_v_0_MPORT_172_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_7_tile_v_3_MPORT_4_en = handshaked & _GEN_1331;
  assign rf_matrix_b_7_tile_v_3_MPORT_4_addr = 8'h43;
  assign rf_matrix_b_7_tile_v_3_MPORT_4_data = rf[rf_matrix_b_7_tile_v_3_MPORT_4_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_7_tile_v_2_MPORT_4_en = handshaked & _GEN_1331;
  assign rf_matrix_b_7_tile_v_2_MPORT_4_addr = 8'h47;
  assign rf_matrix_b_7_tile_v_2_MPORT_4_data = rf[rf_matrix_b_7_tile_v_2_MPORT_4_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_7_tile_v_1_MPORT_4_en = handshaked & _GEN_1331;
  assign rf_matrix_b_7_tile_v_1_MPORT_4_addr = 8'h4b;
  assign rf_matrix_b_7_tile_v_1_MPORT_4_data = rf[rf_matrix_b_7_tile_v_1_MPORT_4_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_7_tile_v_0_MPORT_4_en = handshaked & _GEN_1331;
  assign rf_matrix_b_7_tile_v_0_MPORT_4_addr = 8'h4f;
  assign rf_matrix_b_7_tile_v_0_MPORT_4_data = rf[rf_matrix_b_7_tile_v_0_MPORT_4_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_7_tile_v_3_MPORT_4_en = handshaked & _GEN_1331;
  assign rf_matrix_c_7_tile_v_3_MPORT_4_addr = 8'he6;
  assign rf_matrix_c_7_tile_v_3_MPORT_4_data = rf[rf_matrix_c_7_tile_v_3_MPORT_4_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_7_tile_v_2_MPORT_4_en = handshaked & _GEN_1331;
  assign rf_matrix_c_7_tile_v_2_MPORT_4_addr = 8'he7;
  assign rf_matrix_c_7_tile_v_2_MPORT_4_data = rf[rf_matrix_c_7_tile_v_2_MPORT_4_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_7_tile_v_1_MPORT_4_en = handshaked & _GEN_1331;
  assign rf_matrix_c_7_tile_v_1_MPORT_4_addr = 8'hee;
  assign rf_matrix_c_7_tile_v_1_MPORT_4_data = rf[rf_matrix_c_7_tile_v_1_MPORT_4_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_7_tile_v_0_MPORT_4_en = handshaked & _GEN_1331;
  assign rf_matrix_c_7_tile_v_0_MPORT_4_addr = 8'hef;
  assign rf_matrix_c_7_tile_v_0_MPORT_4_data = rf[rf_matrix_c_7_tile_v_0_MPORT_4_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_1_MPORT_173_en = handshaked & _GEN_1343;
  assign rf_a_tile_v_1_MPORT_173_addr = 8'h38;
  assign rf_a_tile_v_1_MPORT_173_data = rf[rf_a_tile_v_1_MPORT_173_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_0_MPORT_173_en = handshaked & _GEN_1343;
  assign rf_a_tile_v_0_MPORT_173_addr = 8'h3c;
  assign rf_a_tile_v_0_MPORT_173_data = rf[rf_a_tile_v_0_MPORT_173_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_7_tile_v_3_MPORT_5_en = handshaked & _GEN_1343;
  assign rf_matrix_b_7_tile_v_3_MPORT_5_addr = 8'h43;
  assign rf_matrix_b_7_tile_v_3_MPORT_5_data = rf[rf_matrix_b_7_tile_v_3_MPORT_5_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_7_tile_v_2_MPORT_5_en = handshaked & _GEN_1343;
  assign rf_matrix_b_7_tile_v_2_MPORT_5_addr = 8'h47;
  assign rf_matrix_b_7_tile_v_2_MPORT_5_data = rf[rf_matrix_b_7_tile_v_2_MPORT_5_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_7_tile_v_1_MPORT_5_en = handshaked & _GEN_1343;
  assign rf_matrix_b_7_tile_v_1_MPORT_5_addr = 8'h4b;
  assign rf_matrix_b_7_tile_v_1_MPORT_5_data = rf[rf_matrix_b_7_tile_v_1_MPORT_5_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_7_tile_v_0_MPORT_5_en = handshaked & _GEN_1343;
  assign rf_matrix_b_7_tile_v_0_MPORT_5_addr = 8'h4f;
  assign rf_matrix_b_7_tile_v_0_MPORT_5_data = rf[rf_matrix_b_7_tile_v_0_MPORT_5_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_7_tile_v_3_MPORT_5_en = handshaked & _GEN_1343;
  assign rf_matrix_c_7_tile_v_3_MPORT_5_addr = 8'hf6;
  assign rf_matrix_c_7_tile_v_3_MPORT_5_data = rf[rf_matrix_c_7_tile_v_3_MPORT_5_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_7_tile_v_2_MPORT_5_en = handshaked & _GEN_1343;
  assign rf_matrix_c_7_tile_v_2_MPORT_5_addr = 8'hf7;
  assign rf_matrix_c_7_tile_v_2_MPORT_5_data = rf[rf_matrix_c_7_tile_v_2_MPORT_5_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_7_tile_v_1_MPORT_5_en = handshaked & _GEN_1343;
  assign rf_matrix_c_7_tile_v_1_MPORT_5_addr = 8'hfe;
  assign rf_matrix_c_7_tile_v_1_MPORT_5_data = rf[rf_matrix_c_7_tile_v_1_MPORT_5_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_7_tile_v_0_MPORT_5_en = handshaked & _GEN_1343;
  assign rf_matrix_c_7_tile_v_0_MPORT_5_addr = 8'hff;
  assign rf_matrix_c_7_tile_v_0_MPORT_5_data = rf[rf_matrix_c_7_tile_v_0_MPORT_5_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_1_MPORT_174_en = handshaked & _GEN_1355;
  assign rf_a_tile_v_1_MPORT_174_addr = 8'h31;
  assign rf_a_tile_v_1_MPORT_174_data = rf[rf_a_tile_v_1_MPORT_174_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_0_MPORT_174_en = handshaked & _GEN_1355;
  assign rf_a_tile_v_0_MPORT_174_addr = 8'h35;
  assign rf_a_tile_v_0_MPORT_174_data = rf[rf_a_tile_v_0_MPORT_174_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_7_tile_v_3_MPORT_6_en = handshaked & _GEN_1355;
  assign rf_matrix_b_7_tile_v_3_MPORT_6_addr = 8'h53;
  assign rf_matrix_b_7_tile_v_3_MPORT_6_data = rf[rf_matrix_b_7_tile_v_3_MPORT_6_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_7_tile_v_2_MPORT_6_en = handshaked & _GEN_1355;
  assign rf_matrix_b_7_tile_v_2_MPORT_6_addr = 8'h57;
  assign rf_matrix_b_7_tile_v_2_MPORT_6_data = rf[rf_matrix_b_7_tile_v_2_MPORT_6_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_7_tile_v_1_MPORT_6_en = handshaked & _GEN_1355;
  assign rf_matrix_b_7_tile_v_1_MPORT_6_addr = 8'h5b;
  assign rf_matrix_b_7_tile_v_1_MPORT_6_data = rf[rf_matrix_b_7_tile_v_1_MPORT_6_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_7_tile_v_0_MPORT_6_en = handshaked & _GEN_1355;
  assign rf_matrix_b_7_tile_v_0_MPORT_6_addr = 8'h5f;
  assign rf_matrix_b_7_tile_v_0_MPORT_6_data = rf[rf_matrix_b_7_tile_v_0_MPORT_6_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_7_tile_v_3_MPORT_6_en = handshaked & _GEN_1355;
  assign rf_matrix_c_7_tile_v_3_MPORT_6_addr = 8'he4;
  assign rf_matrix_c_7_tile_v_3_MPORT_6_data = rf[rf_matrix_c_7_tile_v_3_MPORT_6_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_7_tile_v_2_MPORT_6_en = handshaked & _GEN_1355;
  assign rf_matrix_c_7_tile_v_2_MPORT_6_addr = 8'he5;
  assign rf_matrix_c_7_tile_v_2_MPORT_6_data = rf[rf_matrix_c_7_tile_v_2_MPORT_6_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_7_tile_v_1_MPORT_6_en = handshaked & _GEN_1355;
  assign rf_matrix_c_7_tile_v_1_MPORT_6_addr = 8'hec;
  assign rf_matrix_c_7_tile_v_1_MPORT_6_data = rf[rf_matrix_c_7_tile_v_1_MPORT_6_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_7_tile_v_0_MPORT_6_en = handshaked & _GEN_1355;
  assign rf_matrix_c_7_tile_v_0_MPORT_6_addr = 8'hed;
  assign rf_matrix_c_7_tile_v_0_MPORT_6_data = rf[rf_matrix_c_7_tile_v_0_MPORT_6_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_3_MPORT_58_en = handshaked & _GEN_1367;
  assign rf_a_tile_v_3_MPORT_58_addr = 8'h31;
  assign rf_a_tile_v_3_MPORT_58_data = rf[rf_a_tile_v_3_MPORT_58_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_2_MPORT_58_en = handshaked & _GEN_1367;
  assign rf_a_tile_v_2_MPORT_58_addr = 8'h35;
  assign rf_a_tile_v_2_MPORT_58_data = rf[rf_a_tile_v_2_MPORT_58_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_1_MPORT_175_en = handshaked & _GEN_1367;
  assign rf_a_tile_v_1_MPORT_175_addr = 8'h39;
  assign rf_a_tile_v_1_MPORT_175_data = rf[rf_a_tile_v_1_MPORT_175_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_0_MPORT_175_en = handshaked & _GEN_1367;
  assign rf_a_tile_v_0_MPORT_175_addr = 8'h3d;
  assign rf_a_tile_v_0_MPORT_175_data = rf[rf_a_tile_v_0_MPORT_175_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_7_tile_v_3_MPORT_7_en = handshaked & _GEN_1367;
  assign rf_matrix_b_7_tile_v_3_MPORT_7_addr = 8'h53;
  assign rf_matrix_b_7_tile_v_3_MPORT_7_data = rf[rf_matrix_b_7_tile_v_3_MPORT_7_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_7_tile_v_2_MPORT_7_en = handshaked & _GEN_1367;
  assign rf_matrix_b_7_tile_v_2_MPORT_7_addr = 8'h57;
  assign rf_matrix_b_7_tile_v_2_MPORT_7_data = rf[rf_matrix_b_7_tile_v_2_MPORT_7_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_7_tile_v_1_MPORT_7_en = handshaked & _GEN_1367;
  assign rf_matrix_b_7_tile_v_1_MPORT_7_addr = 8'h5b;
  assign rf_matrix_b_7_tile_v_1_MPORT_7_data = rf[rf_matrix_b_7_tile_v_1_MPORT_7_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_7_tile_v_0_MPORT_7_en = handshaked & _GEN_1367;
  assign rf_matrix_b_7_tile_v_0_MPORT_7_addr = 8'h5f;
  assign rf_matrix_b_7_tile_v_0_MPORT_7_data = rf[rf_matrix_b_7_tile_v_0_MPORT_7_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_7_tile_v_3_MPORT_7_en = handshaked & _GEN_1367;
  assign rf_matrix_c_7_tile_v_3_MPORT_7_addr = 8'hb2;
  assign rf_matrix_c_7_tile_v_3_MPORT_7_data = rf[rf_matrix_c_7_tile_v_3_MPORT_7_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_7_tile_v_2_MPORT_7_en = handshaked & _GEN_1367;
  assign rf_matrix_c_7_tile_v_2_MPORT_7_addr = 8'hb6;
  assign rf_matrix_c_7_tile_v_2_MPORT_7_data = rf[rf_matrix_c_7_tile_v_2_MPORT_7_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_7_tile_v_1_MPORT_7_en = handshaked & _GEN_1367;
  assign rf_matrix_c_7_tile_v_1_MPORT_7_addr = 8'hba;
  assign rf_matrix_c_7_tile_v_1_MPORT_7_data = rf[rf_matrix_c_7_tile_v_1_MPORT_7_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_7_tile_v_0_MPORT_7_en = handshaked & _GEN_1367;
  assign rf_matrix_c_7_tile_v_0_MPORT_7_addr = 8'hbe;
  assign rf_matrix_c_7_tile_v_0_MPORT_7_data = rf[rf_matrix_c_7_tile_v_0_MPORT_7_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_1_MPORT_176_en = handshaked & _GEN_1381;
  assign rf_a_tile_v_1_MPORT_176_addr = 8'h39;
  assign rf_a_tile_v_1_MPORT_176_data = rf[rf_a_tile_v_1_MPORT_176_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_0_MPORT_176_en = handshaked & _GEN_1381;
  assign rf_a_tile_v_0_MPORT_176_addr = 8'h3d;
  assign rf_a_tile_v_0_MPORT_176_data = rf[rf_a_tile_v_0_MPORT_176_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_7_tile_v_3_MPORT_8_en = handshaked & _GEN_1381;
  assign rf_matrix_b_7_tile_v_3_MPORT_8_addr = 8'h53;
  assign rf_matrix_b_7_tile_v_3_MPORT_8_data = rf[rf_matrix_b_7_tile_v_3_MPORT_8_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_7_tile_v_2_MPORT_8_en = handshaked & _GEN_1381;
  assign rf_matrix_b_7_tile_v_2_MPORT_8_addr = 8'h57;
  assign rf_matrix_b_7_tile_v_2_MPORT_8_data = rf[rf_matrix_b_7_tile_v_2_MPORT_8_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_7_tile_v_1_MPORT_8_en = handshaked & _GEN_1381;
  assign rf_matrix_b_7_tile_v_1_MPORT_8_addr = 8'h5b;
  assign rf_matrix_b_7_tile_v_1_MPORT_8_data = rf[rf_matrix_b_7_tile_v_1_MPORT_8_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_7_tile_v_0_MPORT_8_en = handshaked & _GEN_1381;
  assign rf_matrix_b_7_tile_v_0_MPORT_8_addr = 8'h5f;
  assign rf_matrix_b_7_tile_v_0_MPORT_8_data = rf[rf_matrix_b_7_tile_v_0_MPORT_8_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_7_tile_v_3_MPORT_8_en = handshaked & _GEN_1381;
  assign rf_matrix_c_7_tile_v_3_MPORT_8_addr = 8'hf4;
  assign rf_matrix_c_7_tile_v_3_MPORT_8_data = rf[rf_matrix_c_7_tile_v_3_MPORT_8_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_7_tile_v_2_MPORT_8_en = handshaked & _GEN_1381;
  assign rf_matrix_c_7_tile_v_2_MPORT_8_addr = 8'hf5;
  assign rf_matrix_c_7_tile_v_2_MPORT_8_data = rf[rf_matrix_c_7_tile_v_2_MPORT_8_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_7_tile_v_1_MPORT_8_en = handshaked & _GEN_1381;
  assign rf_matrix_c_7_tile_v_1_MPORT_8_addr = 8'hfc;
  assign rf_matrix_c_7_tile_v_1_MPORT_8_data = rf[rf_matrix_c_7_tile_v_1_MPORT_8_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_7_tile_v_0_MPORT_8_en = handshaked & _GEN_1381;
  assign rf_matrix_c_7_tile_v_0_MPORT_8_addr = 8'hfd;
  assign rf_matrix_c_7_tile_v_0_MPORT_8_data = rf[rf_matrix_c_7_tile_v_0_MPORT_8_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_3_MPORT_59_en = handshaked & _GEN_1393;
  assign rf_a_tile_v_3_MPORT_59_addr = 8'h31;
  assign rf_a_tile_v_3_MPORT_59_data = rf[rf_a_tile_v_3_MPORT_59_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_2_MPORT_59_en = handshaked & _GEN_1393;
  assign rf_a_tile_v_2_MPORT_59_addr = 8'h35;
  assign rf_a_tile_v_2_MPORT_59_data = rf[rf_a_tile_v_2_MPORT_59_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_1_MPORT_177_en = handshaked & _GEN_1393;
  assign rf_a_tile_v_1_MPORT_177_addr = 8'h39;
  assign rf_a_tile_v_1_MPORT_177_data = rf[rf_a_tile_v_1_MPORT_177_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_0_MPORT_177_en = handshaked & _GEN_1393;
  assign rf_a_tile_v_0_MPORT_177_addr = 8'h3d;
  assign rf_a_tile_v_0_MPORT_177_data = rf[rf_a_tile_v_0_MPORT_177_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_7_tile_v_3_MPORT_9_en = handshaked & _GEN_1393;
  assign rf_matrix_b_7_tile_v_3_MPORT_9_addr = 8'h53;
  assign rf_matrix_b_7_tile_v_3_MPORT_9_data = rf[rf_matrix_b_7_tile_v_3_MPORT_9_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_7_tile_v_2_MPORT_9_en = handshaked & _GEN_1393;
  assign rf_matrix_b_7_tile_v_2_MPORT_9_addr = 8'h57;
  assign rf_matrix_b_7_tile_v_2_MPORT_9_data = rf[rf_matrix_b_7_tile_v_2_MPORT_9_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_7_tile_v_1_MPORT_9_en = handshaked & _GEN_1393;
  assign rf_matrix_b_7_tile_v_1_MPORT_9_addr = 8'h5b;
  assign rf_matrix_b_7_tile_v_1_MPORT_9_data = rf[rf_matrix_b_7_tile_v_1_MPORT_9_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_7_tile_v_0_MPORT_9_en = handshaked & _GEN_1393;
  assign rf_matrix_b_7_tile_v_0_MPORT_9_addr = 8'h5f;
  assign rf_matrix_b_7_tile_v_0_MPORT_9_data = rf[rf_matrix_b_7_tile_v_0_MPORT_9_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_7_tile_v_3_MPORT_9_en = handshaked & _GEN_1393;
  assign rf_matrix_c_7_tile_v_3_MPORT_9_addr = 8'hb3;
  assign rf_matrix_c_7_tile_v_3_MPORT_9_data = rf[rf_matrix_c_7_tile_v_3_MPORT_9_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_7_tile_v_2_MPORT_9_en = handshaked & _GEN_1393;
  assign rf_matrix_c_7_tile_v_2_MPORT_9_addr = 8'hb7;
  assign rf_matrix_c_7_tile_v_2_MPORT_9_data = rf[rf_matrix_c_7_tile_v_2_MPORT_9_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_7_tile_v_1_MPORT_9_en = handshaked & _GEN_1393;
  assign rf_matrix_c_7_tile_v_1_MPORT_9_addr = 8'hbb;
  assign rf_matrix_c_7_tile_v_1_MPORT_9_data = rf[rf_matrix_c_7_tile_v_1_MPORT_9_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_7_tile_v_0_MPORT_9_en = handshaked & _GEN_1393;
  assign rf_matrix_c_7_tile_v_0_MPORT_9_addr = 8'hbf;
  assign rf_matrix_c_7_tile_v_0_MPORT_9_data = rf[rf_matrix_c_7_tile_v_0_MPORT_9_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_1_MPORT_178_en = handshaked & _GEN_1407;
  assign rf_a_tile_v_1_MPORT_178_addr = 8'h31;
  assign rf_a_tile_v_1_MPORT_178_data = rf[rf_a_tile_v_1_MPORT_178_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_0_MPORT_178_en = handshaked & _GEN_1407;
  assign rf_a_tile_v_0_MPORT_178_addr = 8'h35;
  assign rf_a_tile_v_0_MPORT_178_data = rf[rf_a_tile_v_0_MPORT_178_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_7_tile_v_3_MPORT_10_en = handshaked & _GEN_1407;
  assign rf_matrix_b_7_tile_v_3_MPORT_10_addr = 8'h53;
  assign rf_matrix_b_7_tile_v_3_MPORT_10_data = rf[rf_matrix_b_7_tile_v_3_MPORT_10_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_7_tile_v_2_MPORT_10_en = handshaked & _GEN_1407;
  assign rf_matrix_b_7_tile_v_2_MPORT_10_addr = 8'h57;
  assign rf_matrix_b_7_tile_v_2_MPORT_10_data = rf[rf_matrix_b_7_tile_v_2_MPORT_10_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_7_tile_v_1_MPORT_10_en = handshaked & _GEN_1407;
  assign rf_matrix_b_7_tile_v_1_MPORT_10_addr = 8'h5b;
  assign rf_matrix_b_7_tile_v_1_MPORT_10_data = rf[rf_matrix_b_7_tile_v_1_MPORT_10_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_7_tile_v_0_MPORT_10_en = handshaked & _GEN_1407;
  assign rf_matrix_b_7_tile_v_0_MPORT_10_addr = 8'h5f;
  assign rf_matrix_b_7_tile_v_0_MPORT_10_data = rf[rf_matrix_b_7_tile_v_0_MPORT_10_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_7_tile_v_3_MPORT_10_en = handshaked & _GEN_1407;
  assign rf_matrix_c_7_tile_v_3_MPORT_10_addr = 8'he6;
  assign rf_matrix_c_7_tile_v_3_MPORT_10_data = rf[rf_matrix_c_7_tile_v_3_MPORT_10_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_7_tile_v_2_MPORT_10_en = handshaked & _GEN_1407;
  assign rf_matrix_c_7_tile_v_2_MPORT_10_addr = 8'he7;
  assign rf_matrix_c_7_tile_v_2_MPORT_10_data = rf[rf_matrix_c_7_tile_v_2_MPORT_10_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_7_tile_v_1_MPORT_10_en = handshaked & _GEN_1407;
  assign rf_matrix_c_7_tile_v_1_MPORT_10_addr = 8'hee;
  assign rf_matrix_c_7_tile_v_1_MPORT_10_data = rf[rf_matrix_c_7_tile_v_1_MPORT_10_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_7_tile_v_0_MPORT_10_en = handshaked & _GEN_1407;
  assign rf_matrix_c_7_tile_v_0_MPORT_10_addr = 8'hef;
  assign rf_matrix_c_7_tile_v_0_MPORT_10_data = rf[rf_matrix_c_7_tile_v_0_MPORT_10_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_1_MPORT_179_en = handshaked & _GEN_1419;
  assign rf_a_tile_v_1_MPORT_179_addr = 8'h39;
  assign rf_a_tile_v_1_MPORT_179_data = rf[rf_a_tile_v_1_MPORT_179_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_0_MPORT_179_en = handshaked & _GEN_1419;
  assign rf_a_tile_v_0_MPORT_179_addr = 8'h3d;
  assign rf_a_tile_v_0_MPORT_179_data = rf[rf_a_tile_v_0_MPORT_179_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_7_tile_v_3_MPORT_11_en = handshaked & _GEN_1419;
  assign rf_matrix_b_7_tile_v_3_MPORT_11_addr = 8'h53;
  assign rf_matrix_b_7_tile_v_3_MPORT_11_data = rf[rf_matrix_b_7_tile_v_3_MPORT_11_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_7_tile_v_2_MPORT_11_en = handshaked & _GEN_1419;
  assign rf_matrix_b_7_tile_v_2_MPORT_11_addr = 8'h57;
  assign rf_matrix_b_7_tile_v_2_MPORT_11_data = rf[rf_matrix_b_7_tile_v_2_MPORT_11_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_7_tile_v_1_MPORT_11_en = handshaked & _GEN_1419;
  assign rf_matrix_b_7_tile_v_1_MPORT_11_addr = 8'h5b;
  assign rf_matrix_b_7_tile_v_1_MPORT_11_data = rf[rf_matrix_b_7_tile_v_1_MPORT_11_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_7_tile_v_0_MPORT_11_en = handshaked & _GEN_1419;
  assign rf_matrix_b_7_tile_v_0_MPORT_11_addr = 8'h5f;
  assign rf_matrix_b_7_tile_v_0_MPORT_11_data = rf[rf_matrix_b_7_tile_v_0_MPORT_11_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_7_tile_v_3_MPORT_11_en = handshaked & _GEN_1419;
  assign rf_matrix_c_7_tile_v_3_MPORT_11_addr = 8'hf6;
  assign rf_matrix_c_7_tile_v_3_MPORT_11_data = rf[rf_matrix_c_7_tile_v_3_MPORT_11_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_7_tile_v_2_MPORT_11_en = handshaked & _GEN_1419;
  assign rf_matrix_c_7_tile_v_2_MPORT_11_addr = 8'hf7;
  assign rf_matrix_c_7_tile_v_2_MPORT_11_data = rf[rf_matrix_c_7_tile_v_2_MPORT_11_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_7_tile_v_1_MPORT_11_en = handshaked & _GEN_1419;
  assign rf_matrix_c_7_tile_v_1_MPORT_11_addr = 8'hfe;
  assign rf_matrix_c_7_tile_v_1_MPORT_11_data = rf[rf_matrix_c_7_tile_v_1_MPORT_11_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_7_tile_v_0_MPORT_11_en = handshaked & _GEN_1419;
  assign rf_matrix_c_7_tile_v_0_MPORT_11_addr = 8'hff;
  assign rf_matrix_c_7_tile_v_0_MPORT_11_data = rf[rf_matrix_c_7_tile_v_0_MPORT_11_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_1_MPORT_180_en = handshaked & _GEN_1431;
  assign rf_a_tile_v_1_MPORT_180_addr = 8'h32;
  assign rf_a_tile_v_1_MPORT_180_data = rf[rf_a_tile_v_1_MPORT_180_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_0_MPORT_180_en = handshaked & _GEN_1431;
  assign rf_a_tile_v_0_MPORT_180_addr = 8'h36;
  assign rf_a_tile_v_0_MPORT_180_data = rf[rf_a_tile_v_0_MPORT_180_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_7_tile_v_3_MPORT_12_en = handshaked & _GEN_1431;
  assign rf_matrix_b_7_tile_v_3_MPORT_12_addr = 8'h63;
  assign rf_matrix_b_7_tile_v_3_MPORT_12_data = rf[rf_matrix_b_7_tile_v_3_MPORT_12_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_7_tile_v_2_MPORT_12_en = handshaked & _GEN_1431;
  assign rf_matrix_b_7_tile_v_2_MPORT_12_addr = 8'h67;
  assign rf_matrix_b_7_tile_v_2_MPORT_12_data = rf[rf_matrix_b_7_tile_v_2_MPORT_12_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_7_tile_v_1_MPORT_12_en = handshaked & _GEN_1431;
  assign rf_matrix_b_7_tile_v_1_MPORT_12_addr = 8'h6b;
  assign rf_matrix_b_7_tile_v_1_MPORT_12_data = rf[rf_matrix_b_7_tile_v_1_MPORT_12_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_7_tile_v_0_MPORT_12_en = handshaked & _GEN_1431;
  assign rf_matrix_b_7_tile_v_0_MPORT_12_addr = 8'h6f;
  assign rf_matrix_b_7_tile_v_0_MPORT_12_data = rf[rf_matrix_b_7_tile_v_0_MPORT_12_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_7_tile_v_3_MPORT_12_en = handshaked & _GEN_1431;
  assign rf_matrix_c_7_tile_v_3_MPORT_12_addr = 8'he4;
  assign rf_matrix_c_7_tile_v_3_MPORT_12_data = rf[rf_matrix_c_7_tile_v_3_MPORT_12_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_7_tile_v_2_MPORT_12_en = handshaked & _GEN_1431;
  assign rf_matrix_c_7_tile_v_2_MPORT_12_addr = 8'he5;
  assign rf_matrix_c_7_tile_v_2_MPORT_12_data = rf[rf_matrix_c_7_tile_v_2_MPORT_12_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_7_tile_v_1_MPORT_12_en = handshaked & _GEN_1431;
  assign rf_matrix_c_7_tile_v_1_MPORT_12_addr = 8'hec;
  assign rf_matrix_c_7_tile_v_1_MPORT_12_data = rf[rf_matrix_c_7_tile_v_1_MPORT_12_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_7_tile_v_0_MPORT_12_en = handshaked & _GEN_1431;
  assign rf_matrix_c_7_tile_v_0_MPORT_12_addr = 8'hed;
  assign rf_matrix_c_7_tile_v_0_MPORT_12_data = rf[rf_matrix_c_7_tile_v_0_MPORT_12_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_3_MPORT_60_en = handshaked & _GEN_1443;
  assign rf_a_tile_v_3_MPORT_60_addr = 8'h32;
  assign rf_a_tile_v_3_MPORT_60_data = rf[rf_a_tile_v_3_MPORT_60_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_2_MPORT_60_en = handshaked & _GEN_1443;
  assign rf_a_tile_v_2_MPORT_60_addr = 8'h36;
  assign rf_a_tile_v_2_MPORT_60_data = rf[rf_a_tile_v_2_MPORT_60_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_1_MPORT_181_en = handshaked & _GEN_1443;
  assign rf_a_tile_v_1_MPORT_181_addr = 8'h3a;
  assign rf_a_tile_v_1_MPORT_181_data = rf[rf_a_tile_v_1_MPORT_181_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_0_MPORT_181_en = handshaked & _GEN_1443;
  assign rf_a_tile_v_0_MPORT_181_addr = 8'h3e;
  assign rf_a_tile_v_0_MPORT_181_data = rf[rf_a_tile_v_0_MPORT_181_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_7_tile_v_3_MPORT_13_en = handshaked & _GEN_1443;
  assign rf_matrix_b_7_tile_v_3_MPORT_13_addr = 8'h63;
  assign rf_matrix_b_7_tile_v_3_MPORT_13_data = rf[rf_matrix_b_7_tile_v_3_MPORT_13_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_7_tile_v_2_MPORT_13_en = handshaked & _GEN_1443;
  assign rf_matrix_b_7_tile_v_2_MPORT_13_addr = 8'h67;
  assign rf_matrix_b_7_tile_v_2_MPORT_13_data = rf[rf_matrix_b_7_tile_v_2_MPORT_13_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_7_tile_v_1_MPORT_13_en = handshaked & _GEN_1443;
  assign rf_matrix_b_7_tile_v_1_MPORT_13_addr = 8'h6b;
  assign rf_matrix_b_7_tile_v_1_MPORT_13_data = rf[rf_matrix_b_7_tile_v_1_MPORT_13_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_7_tile_v_0_MPORT_13_en = handshaked & _GEN_1443;
  assign rf_matrix_b_7_tile_v_0_MPORT_13_addr = 8'h6f;
  assign rf_matrix_b_7_tile_v_0_MPORT_13_data = rf[rf_matrix_b_7_tile_v_0_MPORT_13_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_7_tile_v_3_MPORT_13_en = handshaked & _GEN_1443;
  assign rf_matrix_c_7_tile_v_3_MPORT_13_addr = 8'hb2;
  assign rf_matrix_c_7_tile_v_3_MPORT_13_data = rf[rf_matrix_c_7_tile_v_3_MPORT_13_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_7_tile_v_2_MPORT_13_en = handshaked & _GEN_1443;
  assign rf_matrix_c_7_tile_v_2_MPORT_13_addr = 8'hb6;
  assign rf_matrix_c_7_tile_v_2_MPORT_13_data = rf[rf_matrix_c_7_tile_v_2_MPORT_13_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_7_tile_v_1_MPORT_13_en = handshaked & _GEN_1443;
  assign rf_matrix_c_7_tile_v_1_MPORT_13_addr = 8'hba;
  assign rf_matrix_c_7_tile_v_1_MPORT_13_data = rf[rf_matrix_c_7_tile_v_1_MPORT_13_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_7_tile_v_0_MPORT_13_en = handshaked & _GEN_1443;
  assign rf_matrix_c_7_tile_v_0_MPORT_13_addr = 8'hbe;
  assign rf_matrix_c_7_tile_v_0_MPORT_13_data = rf[rf_matrix_c_7_tile_v_0_MPORT_13_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_1_MPORT_182_en = handshaked & _GEN_1457;
  assign rf_a_tile_v_1_MPORT_182_addr = 8'h3a;
  assign rf_a_tile_v_1_MPORT_182_data = rf[rf_a_tile_v_1_MPORT_182_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_0_MPORT_182_en = handshaked & _GEN_1457;
  assign rf_a_tile_v_0_MPORT_182_addr = 8'h3e;
  assign rf_a_tile_v_0_MPORT_182_data = rf[rf_a_tile_v_0_MPORT_182_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_7_tile_v_3_MPORT_14_en = handshaked & _GEN_1457;
  assign rf_matrix_b_7_tile_v_3_MPORT_14_addr = 8'h63;
  assign rf_matrix_b_7_tile_v_3_MPORT_14_data = rf[rf_matrix_b_7_tile_v_3_MPORT_14_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_7_tile_v_2_MPORT_14_en = handshaked & _GEN_1457;
  assign rf_matrix_b_7_tile_v_2_MPORT_14_addr = 8'h67;
  assign rf_matrix_b_7_tile_v_2_MPORT_14_data = rf[rf_matrix_b_7_tile_v_2_MPORT_14_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_7_tile_v_1_MPORT_14_en = handshaked & _GEN_1457;
  assign rf_matrix_b_7_tile_v_1_MPORT_14_addr = 8'h6b;
  assign rf_matrix_b_7_tile_v_1_MPORT_14_data = rf[rf_matrix_b_7_tile_v_1_MPORT_14_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_7_tile_v_0_MPORT_14_en = handshaked & _GEN_1457;
  assign rf_matrix_b_7_tile_v_0_MPORT_14_addr = 8'h6f;
  assign rf_matrix_b_7_tile_v_0_MPORT_14_data = rf[rf_matrix_b_7_tile_v_0_MPORT_14_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_7_tile_v_3_MPORT_14_en = handshaked & _GEN_1457;
  assign rf_matrix_c_7_tile_v_3_MPORT_14_addr = 8'hf4;
  assign rf_matrix_c_7_tile_v_3_MPORT_14_data = rf[rf_matrix_c_7_tile_v_3_MPORT_14_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_7_tile_v_2_MPORT_14_en = handshaked & _GEN_1457;
  assign rf_matrix_c_7_tile_v_2_MPORT_14_addr = 8'hf5;
  assign rf_matrix_c_7_tile_v_2_MPORT_14_data = rf[rf_matrix_c_7_tile_v_2_MPORT_14_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_7_tile_v_1_MPORT_14_en = handshaked & _GEN_1457;
  assign rf_matrix_c_7_tile_v_1_MPORT_14_addr = 8'hfc;
  assign rf_matrix_c_7_tile_v_1_MPORT_14_data = rf[rf_matrix_c_7_tile_v_1_MPORT_14_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_7_tile_v_0_MPORT_14_en = handshaked & _GEN_1457;
  assign rf_matrix_c_7_tile_v_0_MPORT_14_addr = 8'hfd;
  assign rf_matrix_c_7_tile_v_0_MPORT_14_data = rf[rf_matrix_c_7_tile_v_0_MPORT_14_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_3_MPORT_61_en = handshaked & _GEN_1469;
  assign rf_a_tile_v_3_MPORT_61_addr = 8'h32;
  assign rf_a_tile_v_3_MPORT_61_data = rf[rf_a_tile_v_3_MPORT_61_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_2_MPORT_61_en = handshaked & _GEN_1469;
  assign rf_a_tile_v_2_MPORT_61_addr = 8'h36;
  assign rf_a_tile_v_2_MPORT_61_data = rf[rf_a_tile_v_2_MPORT_61_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_1_MPORT_183_en = handshaked & _GEN_1469;
  assign rf_a_tile_v_1_MPORT_183_addr = 8'h3a;
  assign rf_a_tile_v_1_MPORT_183_data = rf[rf_a_tile_v_1_MPORT_183_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_0_MPORT_183_en = handshaked & _GEN_1469;
  assign rf_a_tile_v_0_MPORT_183_addr = 8'h3e;
  assign rf_a_tile_v_0_MPORT_183_data = rf[rf_a_tile_v_0_MPORT_183_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_7_tile_v_3_MPORT_15_en = handshaked & _GEN_1469;
  assign rf_matrix_b_7_tile_v_3_MPORT_15_addr = 8'h63;
  assign rf_matrix_b_7_tile_v_3_MPORT_15_data = rf[rf_matrix_b_7_tile_v_3_MPORT_15_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_7_tile_v_2_MPORT_15_en = handshaked & _GEN_1469;
  assign rf_matrix_b_7_tile_v_2_MPORT_15_addr = 8'h67;
  assign rf_matrix_b_7_tile_v_2_MPORT_15_data = rf[rf_matrix_b_7_tile_v_2_MPORT_15_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_7_tile_v_1_MPORT_15_en = handshaked & _GEN_1469;
  assign rf_matrix_b_7_tile_v_1_MPORT_15_addr = 8'h6b;
  assign rf_matrix_b_7_tile_v_1_MPORT_15_data = rf[rf_matrix_b_7_tile_v_1_MPORT_15_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_7_tile_v_0_MPORT_15_en = handshaked & _GEN_1469;
  assign rf_matrix_b_7_tile_v_0_MPORT_15_addr = 8'h6f;
  assign rf_matrix_b_7_tile_v_0_MPORT_15_data = rf[rf_matrix_b_7_tile_v_0_MPORT_15_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_7_tile_v_3_MPORT_15_en = handshaked & _GEN_1469;
  assign rf_matrix_c_7_tile_v_3_MPORT_15_addr = 8'hb3;
  assign rf_matrix_c_7_tile_v_3_MPORT_15_data = rf[rf_matrix_c_7_tile_v_3_MPORT_15_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_7_tile_v_2_MPORT_15_en = handshaked & _GEN_1469;
  assign rf_matrix_c_7_tile_v_2_MPORT_15_addr = 8'hb7;
  assign rf_matrix_c_7_tile_v_2_MPORT_15_data = rf[rf_matrix_c_7_tile_v_2_MPORT_15_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_7_tile_v_1_MPORT_15_en = handshaked & _GEN_1469;
  assign rf_matrix_c_7_tile_v_1_MPORT_15_addr = 8'hbb;
  assign rf_matrix_c_7_tile_v_1_MPORT_15_data = rf[rf_matrix_c_7_tile_v_1_MPORT_15_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_7_tile_v_0_MPORT_15_en = handshaked & _GEN_1469;
  assign rf_matrix_c_7_tile_v_0_MPORT_15_addr = 8'hbf;
  assign rf_matrix_c_7_tile_v_0_MPORT_15_data = rf[rf_matrix_c_7_tile_v_0_MPORT_15_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_1_MPORT_184_en = handshaked & _GEN_1483;
  assign rf_a_tile_v_1_MPORT_184_addr = 8'h32;
  assign rf_a_tile_v_1_MPORT_184_data = rf[rf_a_tile_v_1_MPORT_184_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_0_MPORT_184_en = handshaked & _GEN_1483;
  assign rf_a_tile_v_0_MPORT_184_addr = 8'h36;
  assign rf_a_tile_v_0_MPORT_184_data = rf[rf_a_tile_v_0_MPORT_184_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_7_tile_v_3_MPORT_16_en = handshaked & _GEN_1483;
  assign rf_matrix_b_7_tile_v_3_MPORT_16_addr = 8'h63;
  assign rf_matrix_b_7_tile_v_3_MPORT_16_data = rf[rf_matrix_b_7_tile_v_3_MPORT_16_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_7_tile_v_2_MPORT_16_en = handshaked & _GEN_1483;
  assign rf_matrix_b_7_tile_v_2_MPORT_16_addr = 8'h67;
  assign rf_matrix_b_7_tile_v_2_MPORT_16_data = rf[rf_matrix_b_7_tile_v_2_MPORT_16_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_7_tile_v_1_MPORT_16_en = handshaked & _GEN_1483;
  assign rf_matrix_b_7_tile_v_1_MPORT_16_addr = 8'h6b;
  assign rf_matrix_b_7_tile_v_1_MPORT_16_data = rf[rf_matrix_b_7_tile_v_1_MPORT_16_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_7_tile_v_0_MPORT_16_en = handshaked & _GEN_1483;
  assign rf_matrix_b_7_tile_v_0_MPORT_16_addr = 8'h6f;
  assign rf_matrix_b_7_tile_v_0_MPORT_16_data = rf[rf_matrix_b_7_tile_v_0_MPORT_16_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_7_tile_v_3_MPORT_16_en = handshaked & _GEN_1483;
  assign rf_matrix_c_7_tile_v_3_MPORT_16_addr = 8'he6;
  assign rf_matrix_c_7_tile_v_3_MPORT_16_data = rf[rf_matrix_c_7_tile_v_3_MPORT_16_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_7_tile_v_2_MPORT_16_en = handshaked & _GEN_1483;
  assign rf_matrix_c_7_tile_v_2_MPORT_16_addr = 8'he7;
  assign rf_matrix_c_7_tile_v_2_MPORT_16_data = rf[rf_matrix_c_7_tile_v_2_MPORT_16_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_7_tile_v_1_MPORT_16_en = handshaked & _GEN_1483;
  assign rf_matrix_c_7_tile_v_1_MPORT_16_addr = 8'hee;
  assign rf_matrix_c_7_tile_v_1_MPORT_16_data = rf[rf_matrix_c_7_tile_v_1_MPORT_16_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_7_tile_v_0_MPORT_16_en = handshaked & _GEN_1483;
  assign rf_matrix_c_7_tile_v_0_MPORT_16_addr = 8'hef;
  assign rf_matrix_c_7_tile_v_0_MPORT_16_data = rf[rf_matrix_c_7_tile_v_0_MPORT_16_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_1_MPORT_185_en = handshaked & _GEN_1495;
  assign rf_a_tile_v_1_MPORT_185_addr = 8'h3a;
  assign rf_a_tile_v_1_MPORT_185_data = rf[rf_a_tile_v_1_MPORT_185_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_0_MPORT_185_en = handshaked & _GEN_1495;
  assign rf_a_tile_v_0_MPORT_185_addr = 8'h3e;
  assign rf_a_tile_v_0_MPORT_185_data = rf[rf_a_tile_v_0_MPORT_185_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_7_tile_v_3_MPORT_17_en = handshaked & _GEN_1495;
  assign rf_matrix_b_7_tile_v_3_MPORT_17_addr = 8'h63;
  assign rf_matrix_b_7_tile_v_3_MPORT_17_data = rf[rf_matrix_b_7_tile_v_3_MPORT_17_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_7_tile_v_2_MPORT_17_en = handshaked & _GEN_1495;
  assign rf_matrix_b_7_tile_v_2_MPORT_17_addr = 8'h67;
  assign rf_matrix_b_7_tile_v_2_MPORT_17_data = rf[rf_matrix_b_7_tile_v_2_MPORT_17_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_7_tile_v_1_MPORT_17_en = handshaked & _GEN_1495;
  assign rf_matrix_b_7_tile_v_1_MPORT_17_addr = 8'h6b;
  assign rf_matrix_b_7_tile_v_1_MPORT_17_data = rf[rf_matrix_b_7_tile_v_1_MPORT_17_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_7_tile_v_0_MPORT_17_en = handshaked & _GEN_1495;
  assign rf_matrix_b_7_tile_v_0_MPORT_17_addr = 8'h6f;
  assign rf_matrix_b_7_tile_v_0_MPORT_17_data = rf[rf_matrix_b_7_tile_v_0_MPORT_17_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_7_tile_v_3_MPORT_17_en = handshaked & _GEN_1495;
  assign rf_matrix_c_7_tile_v_3_MPORT_17_addr = 8'hf6;
  assign rf_matrix_c_7_tile_v_3_MPORT_17_data = rf[rf_matrix_c_7_tile_v_3_MPORT_17_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_7_tile_v_2_MPORT_17_en = handshaked & _GEN_1495;
  assign rf_matrix_c_7_tile_v_2_MPORT_17_addr = 8'hf7;
  assign rf_matrix_c_7_tile_v_2_MPORT_17_data = rf[rf_matrix_c_7_tile_v_2_MPORT_17_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_7_tile_v_1_MPORT_17_en = handshaked & _GEN_1495;
  assign rf_matrix_c_7_tile_v_1_MPORT_17_addr = 8'hfe;
  assign rf_matrix_c_7_tile_v_1_MPORT_17_data = rf[rf_matrix_c_7_tile_v_1_MPORT_17_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_7_tile_v_0_MPORT_17_en = handshaked & _GEN_1495;
  assign rf_matrix_c_7_tile_v_0_MPORT_17_addr = 8'hff;
  assign rf_matrix_c_7_tile_v_0_MPORT_17_data = rf[rf_matrix_c_7_tile_v_0_MPORT_17_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_1_MPORT_186_en = handshaked & _GEN_1507;
  assign rf_a_tile_v_1_MPORT_186_addr = 8'h33;
  assign rf_a_tile_v_1_MPORT_186_data = rf[rf_a_tile_v_1_MPORT_186_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_0_MPORT_186_en = handshaked & _GEN_1507;
  assign rf_a_tile_v_0_MPORT_186_addr = 8'h37;
  assign rf_a_tile_v_0_MPORT_186_data = rf[rf_a_tile_v_0_MPORT_186_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_7_tile_v_3_MPORT_18_en = handshaked & _GEN_1507;
  assign rf_matrix_b_7_tile_v_3_MPORT_18_addr = 8'h73;
  assign rf_matrix_b_7_tile_v_3_MPORT_18_data = rf[rf_matrix_b_7_tile_v_3_MPORT_18_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_7_tile_v_2_MPORT_18_en = handshaked & _GEN_1507;
  assign rf_matrix_b_7_tile_v_2_MPORT_18_addr = 8'h77;
  assign rf_matrix_b_7_tile_v_2_MPORT_18_data = rf[rf_matrix_b_7_tile_v_2_MPORT_18_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_7_tile_v_1_MPORT_18_en = handshaked & _GEN_1507;
  assign rf_matrix_b_7_tile_v_1_MPORT_18_addr = 8'h7b;
  assign rf_matrix_b_7_tile_v_1_MPORT_18_data = rf[rf_matrix_b_7_tile_v_1_MPORT_18_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_7_tile_v_0_MPORT_18_en = handshaked & _GEN_1507;
  assign rf_matrix_b_7_tile_v_0_MPORT_18_addr = 8'h7f;
  assign rf_matrix_b_7_tile_v_0_MPORT_18_data = rf[rf_matrix_b_7_tile_v_0_MPORT_18_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_7_tile_v_3_MPORT_18_en = handshaked & _GEN_1507;
  assign rf_matrix_c_7_tile_v_3_MPORT_18_addr = 8'he4;
  assign rf_matrix_c_7_tile_v_3_MPORT_18_data = rf[rf_matrix_c_7_tile_v_3_MPORT_18_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_7_tile_v_2_MPORT_18_en = handshaked & _GEN_1507;
  assign rf_matrix_c_7_tile_v_2_MPORT_18_addr = 8'he5;
  assign rf_matrix_c_7_tile_v_2_MPORT_18_data = rf[rf_matrix_c_7_tile_v_2_MPORT_18_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_7_tile_v_1_MPORT_18_en = handshaked & _GEN_1507;
  assign rf_matrix_c_7_tile_v_1_MPORT_18_addr = 8'hec;
  assign rf_matrix_c_7_tile_v_1_MPORT_18_data = rf[rf_matrix_c_7_tile_v_1_MPORT_18_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_7_tile_v_0_MPORT_18_en = handshaked & _GEN_1507;
  assign rf_matrix_c_7_tile_v_0_MPORT_18_addr = 8'hed;
  assign rf_matrix_c_7_tile_v_0_MPORT_18_data = rf[rf_matrix_c_7_tile_v_0_MPORT_18_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_3_MPORT_62_en = handshaked & _GEN_1519;
  assign rf_a_tile_v_3_MPORT_62_addr = 8'h33;
  assign rf_a_tile_v_3_MPORT_62_data = rf[rf_a_tile_v_3_MPORT_62_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_2_MPORT_62_en = handshaked & _GEN_1519;
  assign rf_a_tile_v_2_MPORT_62_addr = 8'h37;
  assign rf_a_tile_v_2_MPORT_62_data = rf[rf_a_tile_v_2_MPORT_62_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_1_MPORT_187_en = handshaked & _GEN_1519;
  assign rf_a_tile_v_1_MPORT_187_addr = 8'h3b;
  assign rf_a_tile_v_1_MPORT_187_data = rf[rf_a_tile_v_1_MPORT_187_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_0_MPORT_187_en = handshaked & _GEN_1519;
  assign rf_a_tile_v_0_MPORT_187_addr = 8'h3f;
  assign rf_a_tile_v_0_MPORT_187_data = rf[rf_a_tile_v_0_MPORT_187_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_7_tile_v_3_MPORT_19_en = handshaked & _GEN_1519;
  assign rf_matrix_b_7_tile_v_3_MPORT_19_addr = 8'h73;
  assign rf_matrix_b_7_tile_v_3_MPORT_19_data = rf[rf_matrix_b_7_tile_v_3_MPORT_19_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_7_tile_v_2_MPORT_19_en = handshaked & _GEN_1519;
  assign rf_matrix_b_7_tile_v_2_MPORT_19_addr = 8'h77;
  assign rf_matrix_b_7_tile_v_2_MPORT_19_data = rf[rf_matrix_b_7_tile_v_2_MPORT_19_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_7_tile_v_1_MPORT_19_en = handshaked & _GEN_1519;
  assign rf_matrix_b_7_tile_v_1_MPORT_19_addr = 8'h7b;
  assign rf_matrix_b_7_tile_v_1_MPORT_19_data = rf[rf_matrix_b_7_tile_v_1_MPORT_19_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_7_tile_v_0_MPORT_19_en = handshaked & _GEN_1519;
  assign rf_matrix_b_7_tile_v_0_MPORT_19_addr = 8'h7f;
  assign rf_matrix_b_7_tile_v_0_MPORT_19_data = rf[rf_matrix_b_7_tile_v_0_MPORT_19_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_7_tile_v_3_MPORT_19_en = handshaked & _GEN_1519;
  assign rf_matrix_c_7_tile_v_3_MPORT_19_addr = 8'hb2;
  assign rf_matrix_c_7_tile_v_3_MPORT_19_data = rf[rf_matrix_c_7_tile_v_3_MPORT_19_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_7_tile_v_2_MPORT_19_en = handshaked & _GEN_1519;
  assign rf_matrix_c_7_tile_v_2_MPORT_19_addr = 8'hb6;
  assign rf_matrix_c_7_tile_v_2_MPORT_19_data = rf[rf_matrix_c_7_tile_v_2_MPORT_19_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_7_tile_v_1_MPORT_19_en = handshaked & _GEN_1519;
  assign rf_matrix_c_7_tile_v_1_MPORT_19_addr = 8'hba;
  assign rf_matrix_c_7_tile_v_1_MPORT_19_data = rf[rf_matrix_c_7_tile_v_1_MPORT_19_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_7_tile_v_0_MPORT_19_en = handshaked & _GEN_1519;
  assign rf_matrix_c_7_tile_v_0_MPORT_19_addr = 8'hbe;
  assign rf_matrix_c_7_tile_v_0_MPORT_19_data = rf[rf_matrix_c_7_tile_v_0_MPORT_19_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_1_MPORT_188_en = handshaked & _GEN_1533;
  assign rf_a_tile_v_1_MPORT_188_addr = 8'h3b;
  assign rf_a_tile_v_1_MPORT_188_data = rf[rf_a_tile_v_1_MPORT_188_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_0_MPORT_188_en = handshaked & _GEN_1533;
  assign rf_a_tile_v_0_MPORT_188_addr = 8'h3f;
  assign rf_a_tile_v_0_MPORT_188_data = rf[rf_a_tile_v_0_MPORT_188_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_7_tile_v_3_MPORT_20_en = handshaked & _GEN_1533;
  assign rf_matrix_b_7_tile_v_3_MPORT_20_addr = 8'h73;
  assign rf_matrix_b_7_tile_v_3_MPORT_20_data = rf[rf_matrix_b_7_tile_v_3_MPORT_20_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_7_tile_v_2_MPORT_20_en = handshaked & _GEN_1533;
  assign rf_matrix_b_7_tile_v_2_MPORT_20_addr = 8'h77;
  assign rf_matrix_b_7_tile_v_2_MPORT_20_data = rf[rf_matrix_b_7_tile_v_2_MPORT_20_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_7_tile_v_1_MPORT_20_en = handshaked & _GEN_1533;
  assign rf_matrix_b_7_tile_v_1_MPORT_20_addr = 8'h7b;
  assign rf_matrix_b_7_tile_v_1_MPORT_20_data = rf[rf_matrix_b_7_tile_v_1_MPORT_20_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_7_tile_v_0_MPORT_20_en = handshaked & _GEN_1533;
  assign rf_matrix_b_7_tile_v_0_MPORT_20_addr = 8'h7f;
  assign rf_matrix_b_7_tile_v_0_MPORT_20_data = rf[rf_matrix_b_7_tile_v_0_MPORT_20_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_7_tile_v_3_MPORT_20_en = handshaked & _GEN_1533;
  assign rf_matrix_c_7_tile_v_3_MPORT_20_addr = 8'hf4;
  assign rf_matrix_c_7_tile_v_3_MPORT_20_data = rf[rf_matrix_c_7_tile_v_3_MPORT_20_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_7_tile_v_2_MPORT_20_en = handshaked & _GEN_1533;
  assign rf_matrix_c_7_tile_v_2_MPORT_20_addr = 8'hf5;
  assign rf_matrix_c_7_tile_v_2_MPORT_20_data = rf[rf_matrix_c_7_tile_v_2_MPORT_20_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_7_tile_v_1_MPORT_20_en = handshaked & _GEN_1533;
  assign rf_matrix_c_7_tile_v_1_MPORT_20_addr = 8'hfc;
  assign rf_matrix_c_7_tile_v_1_MPORT_20_data = rf[rf_matrix_c_7_tile_v_1_MPORT_20_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_7_tile_v_0_MPORT_20_en = handshaked & _GEN_1533;
  assign rf_matrix_c_7_tile_v_0_MPORT_20_addr = 8'hfd;
  assign rf_matrix_c_7_tile_v_0_MPORT_20_data = rf[rf_matrix_c_7_tile_v_0_MPORT_20_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_3_MPORT_63_en = handshaked & _GEN_1545;
  assign rf_a_tile_v_3_MPORT_63_addr = 8'h33;
  assign rf_a_tile_v_3_MPORT_63_data = rf[rf_a_tile_v_3_MPORT_63_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_2_MPORT_63_en = handshaked & _GEN_1545;
  assign rf_a_tile_v_2_MPORT_63_addr = 8'h37;
  assign rf_a_tile_v_2_MPORT_63_data = rf[rf_a_tile_v_2_MPORT_63_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_1_MPORT_189_en = handshaked & _GEN_1545;
  assign rf_a_tile_v_1_MPORT_189_addr = 8'h3b;
  assign rf_a_tile_v_1_MPORT_189_data = rf[rf_a_tile_v_1_MPORT_189_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_0_MPORT_189_en = handshaked & _GEN_1545;
  assign rf_a_tile_v_0_MPORT_189_addr = 8'h3f;
  assign rf_a_tile_v_0_MPORT_189_data = rf[rf_a_tile_v_0_MPORT_189_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_7_tile_v_3_MPORT_21_en = handshaked & _GEN_1545;
  assign rf_matrix_b_7_tile_v_3_MPORT_21_addr = 8'h73;
  assign rf_matrix_b_7_tile_v_3_MPORT_21_data = rf[rf_matrix_b_7_tile_v_3_MPORT_21_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_7_tile_v_2_MPORT_21_en = handshaked & _GEN_1545;
  assign rf_matrix_b_7_tile_v_2_MPORT_21_addr = 8'h77;
  assign rf_matrix_b_7_tile_v_2_MPORT_21_data = rf[rf_matrix_b_7_tile_v_2_MPORT_21_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_7_tile_v_1_MPORT_21_en = handshaked & _GEN_1545;
  assign rf_matrix_b_7_tile_v_1_MPORT_21_addr = 8'h7b;
  assign rf_matrix_b_7_tile_v_1_MPORT_21_data = rf[rf_matrix_b_7_tile_v_1_MPORT_21_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_7_tile_v_0_MPORT_21_en = handshaked & _GEN_1545;
  assign rf_matrix_b_7_tile_v_0_MPORT_21_addr = 8'h7f;
  assign rf_matrix_b_7_tile_v_0_MPORT_21_data = rf[rf_matrix_b_7_tile_v_0_MPORT_21_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_7_tile_v_3_MPORT_21_en = handshaked & _GEN_1545;
  assign rf_matrix_c_7_tile_v_3_MPORT_21_addr = 8'hb3;
  assign rf_matrix_c_7_tile_v_3_MPORT_21_data = rf[rf_matrix_c_7_tile_v_3_MPORT_21_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_7_tile_v_2_MPORT_21_en = handshaked & _GEN_1545;
  assign rf_matrix_c_7_tile_v_2_MPORT_21_addr = 8'hb7;
  assign rf_matrix_c_7_tile_v_2_MPORT_21_data = rf[rf_matrix_c_7_tile_v_2_MPORT_21_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_7_tile_v_1_MPORT_21_en = handshaked & _GEN_1545;
  assign rf_matrix_c_7_tile_v_1_MPORT_21_addr = 8'hbb;
  assign rf_matrix_c_7_tile_v_1_MPORT_21_data = rf[rf_matrix_c_7_tile_v_1_MPORT_21_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_7_tile_v_0_MPORT_21_en = handshaked & _GEN_1545;
  assign rf_matrix_c_7_tile_v_0_MPORT_21_addr = 8'hbf;
  assign rf_matrix_c_7_tile_v_0_MPORT_21_data = rf[rf_matrix_c_7_tile_v_0_MPORT_21_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_1_MPORT_190_en = handshaked & _GEN_1559;
  assign rf_a_tile_v_1_MPORT_190_addr = 8'h33;
  assign rf_a_tile_v_1_MPORT_190_data = rf[rf_a_tile_v_1_MPORT_190_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_0_MPORT_190_en = handshaked & _GEN_1559;
  assign rf_a_tile_v_0_MPORT_190_addr = 8'h37;
  assign rf_a_tile_v_0_MPORT_190_data = rf[rf_a_tile_v_0_MPORT_190_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_7_tile_v_3_MPORT_22_en = handshaked & _GEN_1559;
  assign rf_matrix_b_7_tile_v_3_MPORT_22_addr = 8'h73;
  assign rf_matrix_b_7_tile_v_3_MPORT_22_data = rf[rf_matrix_b_7_tile_v_3_MPORT_22_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_7_tile_v_2_MPORT_22_en = handshaked & _GEN_1559;
  assign rf_matrix_b_7_tile_v_2_MPORT_22_addr = 8'h77;
  assign rf_matrix_b_7_tile_v_2_MPORT_22_data = rf[rf_matrix_b_7_tile_v_2_MPORT_22_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_7_tile_v_1_MPORT_22_en = handshaked & _GEN_1559;
  assign rf_matrix_b_7_tile_v_1_MPORT_22_addr = 8'h7b;
  assign rf_matrix_b_7_tile_v_1_MPORT_22_data = rf[rf_matrix_b_7_tile_v_1_MPORT_22_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_7_tile_v_0_MPORT_22_en = handshaked & _GEN_1559;
  assign rf_matrix_b_7_tile_v_0_MPORT_22_addr = 8'h7f;
  assign rf_matrix_b_7_tile_v_0_MPORT_22_data = rf[rf_matrix_b_7_tile_v_0_MPORT_22_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_7_tile_v_3_MPORT_22_en = handshaked & _GEN_1559;
  assign rf_matrix_c_7_tile_v_3_MPORT_22_addr = 8'he6;
  assign rf_matrix_c_7_tile_v_3_MPORT_22_data = rf[rf_matrix_c_7_tile_v_3_MPORT_22_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_7_tile_v_2_MPORT_22_en = handshaked & _GEN_1559;
  assign rf_matrix_c_7_tile_v_2_MPORT_22_addr = 8'he7;
  assign rf_matrix_c_7_tile_v_2_MPORT_22_data = rf[rf_matrix_c_7_tile_v_2_MPORT_22_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_7_tile_v_1_MPORT_22_en = handshaked & _GEN_1559;
  assign rf_matrix_c_7_tile_v_1_MPORT_22_addr = 8'hee;
  assign rf_matrix_c_7_tile_v_1_MPORT_22_data = rf[rf_matrix_c_7_tile_v_1_MPORT_22_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_7_tile_v_0_MPORT_22_en = handshaked & _GEN_1559;
  assign rf_matrix_c_7_tile_v_0_MPORT_22_addr = 8'hef;
  assign rf_matrix_c_7_tile_v_0_MPORT_22_data = rf[rf_matrix_c_7_tile_v_0_MPORT_22_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_1_MPORT_191_en = handshaked & _GEN_1571;
  assign rf_a_tile_v_1_MPORT_191_addr = 8'h3b;
  assign rf_a_tile_v_1_MPORT_191_data = rf[rf_a_tile_v_1_MPORT_191_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_a_tile_v_0_MPORT_191_en = handshaked & _GEN_1571;
  assign rf_a_tile_v_0_MPORT_191_addr = 8'h3f;
  assign rf_a_tile_v_0_MPORT_191_data = rf[rf_a_tile_v_0_MPORT_191_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_7_tile_v_3_MPORT_23_en = handshaked & _GEN_1571;
  assign rf_matrix_b_7_tile_v_3_MPORT_23_addr = 8'h73;
  assign rf_matrix_b_7_tile_v_3_MPORT_23_data = rf[rf_matrix_b_7_tile_v_3_MPORT_23_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_7_tile_v_2_MPORT_23_en = handshaked & _GEN_1571;
  assign rf_matrix_b_7_tile_v_2_MPORT_23_addr = 8'h77;
  assign rf_matrix_b_7_tile_v_2_MPORT_23_data = rf[rf_matrix_b_7_tile_v_2_MPORT_23_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_7_tile_v_1_MPORT_23_en = handshaked & _GEN_1571;
  assign rf_matrix_b_7_tile_v_1_MPORT_23_addr = 8'h7b;
  assign rf_matrix_b_7_tile_v_1_MPORT_23_data = rf[rf_matrix_b_7_tile_v_1_MPORT_23_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_b_7_tile_v_0_MPORT_23_en = handshaked & _GEN_1571;
  assign rf_matrix_b_7_tile_v_0_MPORT_23_addr = 8'h7f;
  assign rf_matrix_b_7_tile_v_0_MPORT_23_data = rf[rf_matrix_b_7_tile_v_0_MPORT_23_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_7_tile_v_3_MPORT_23_en = handshaked & _GEN_1571;
  assign rf_matrix_c_7_tile_v_3_MPORT_23_addr = 8'hf6;
  assign rf_matrix_c_7_tile_v_3_MPORT_23_data = rf[rf_matrix_c_7_tile_v_3_MPORT_23_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_7_tile_v_2_MPORT_23_en = handshaked & _GEN_1571;
  assign rf_matrix_c_7_tile_v_2_MPORT_23_addr = 8'hf7;
  assign rf_matrix_c_7_tile_v_2_MPORT_23_data = rf[rf_matrix_c_7_tile_v_2_MPORT_23_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_7_tile_v_1_MPORT_23_en = handshaked & _GEN_1571;
  assign rf_matrix_c_7_tile_v_1_MPORT_23_addr = 8'hfe;
  assign rf_matrix_c_7_tile_v_1_MPORT_23_data = rf[rf_matrix_c_7_tile_v_1_MPORT_23_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_matrix_c_7_tile_v_0_MPORT_23_en = handshaked & _GEN_1571;
  assign rf_matrix_c_7_tile_v_0_MPORT_23_addr = 8'hff;
  assign rf_matrix_c_7_tile_v_0_MPORT_23_data = rf[rf_matrix_c_7_tile_v_0_MPORT_23_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_io_uart_rf_r_data_MPORT_en = 1'h1;
  assign rf_io_uart_rf_r_data_MPORT_addr = io_uart_rf_r_addr;
  assign rf_io_uart_rf_r_data_MPORT_data = rf[rf_io_uart_rf_r_data_MPORT_addr]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
  assign rf_MPORT_data = io_top_wb_bits_tc0_octet0_threadgroup0_matrix_d_data[255:192];
  assign rf_MPORT_addr = 8'h80;
  assign rf_MPORT_mask = 1'h1;
  assign rf_MPORT_en = _T_162 & _GEN_15391;
  assign rf_MPORT_1_data = io_top_wb_bits_tc0_octet0_threadgroup0_matrix_d_data[191:128];
  assign rf_MPORT_1_addr = 8'h81;
  assign rf_MPORT_1_mask = 1'h1;
  assign rf_MPORT_1_en = _T_162 & _GEN_15391;
  assign rf_MPORT_2_data = io_top_wb_bits_tc0_octet0_threadgroup0_matrix_d_data[127:64];
  assign rf_MPORT_2_addr = 8'h88;
  assign rf_MPORT_2_mask = 1'h1;
  assign rf_MPORT_2_en = _T_162 & _GEN_15391;
  assign rf_MPORT_3_data = io_top_wb_bits_tc0_octet0_threadgroup0_matrix_d_data[63:0];
  assign rf_MPORT_3_addr = 8'h89;
  assign rf_MPORT_3_mask = 1'h1;
  assign rf_MPORT_3_en = _T_162 & _GEN_15391;
  assign rf_MPORT_4_data = io_top_wb_bits_tc0_octet0_threadgroup4_matrix_d_data[255:192];
  assign rf_MPORT_4_addr = 8'ha0;
  assign rf_MPORT_4_mask = 1'h1;
  assign rf_MPORT_4_en = _T_162 & _GEN_15391;
  assign rf_MPORT_5_data = io_top_wb_bits_tc0_octet0_threadgroup4_matrix_d_data[191:128];
  assign rf_MPORT_5_addr = 8'ha1;
  assign rf_MPORT_5_mask = 1'h1;
  assign rf_MPORT_5_en = _T_162 & _GEN_15391;
  assign rf_MPORT_6_data = io_top_wb_bits_tc0_octet0_threadgroup4_matrix_d_data[127:64];
  assign rf_MPORT_6_addr = 8'ha8;
  assign rf_MPORT_6_mask = 1'h1;
  assign rf_MPORT_6_en = _T_162 & _GEN_15391;
  assign rf_MPORT_7_data = io_top_wb_bits_tc0_octet0_threadgroup4_matrix_d_data[63:0];
  assign rf_MPORT_7_addr = 8'ha9;
  assign rf_MPORT_7_mask = 1'h1;
  assign rf_MPORT_7_en = _T_162 & _GEN_15391;
  assign rf_MPORT_8_data = io_top_wb_bits_tc0_octet1_threadgroup0_matrix_d_data[255:192];
  assign rf_MPORT_8_addr = 8'hc0;
  assign rf_MPORT_8_mask = 1'h1;
  assign rf_MPORT_8_en = _T_162 & _GEN_15391;
  assign rf_MPORT_9_data = io_top_wb_bits_tc0_octet1_threadgroup0_matrix_d_data[191:128];
  assign rf_MPORT_9_addr = 8'hc1;
  assign rf_MPORT_9_mask = 1'h1;
  assign rf_MPORT_9_en = _T_162 & _GEN_15391;
  assign rf_MPORT_10_data = io_top_wb_bits_tc0_octet1_threadgroup0_matrix_d_data[127:64];
  assign rf_MPORT_10_addr = 8'hc8;
  assign rf_MPORT_10_mask = 1'h1;
  assign rf_MPORT_10_en = _T_162 & _GEN_15391;
  assign rf_MPORT_11_data = io_top_wb_bits_tc0_octet1_threadgroup0_matrix_d_data[63:0];
  assign rf_MPORT_11_addr = 8'hc9;
  assign rf_MPORT_11_mask = 1'h1;
  assign rf_MPORT_11_en = _T_162 & _GEN_15391;
  assign rf_MPORT_12_data = io_top_wb_bits_tc0_octet1_threadgroup4_matrix_d_data[255:192];
  assign rf_MPORT_12_addr = 8'he0;
  assign rf_MPORT_12_mask = 1'h1;
  assign rf_MPORT_12_en = _T_162 & _GEN_15391;
  assign rf_MPORT_13_data = io_top_wb_bits_tc0_octet1_threadgroup4_matrix_d_data[191:128];
  assign rf_MPORT_13_addr = 8'he1;
  assign rf_MPORT_13_mask = 1'h1;
  assign rf_MPORT_13_en = _T_162 & _GEN_15391;
  assign rf_MPORT_14_data = io_top_wb_bits_tc0_octet1_threadgroup4_matrix_d_data[127:64];
  assign rf_MPORT_14_addr = 8'he8;
  assign rf_MPORT_14_mask = 1'h1;
  assign rf_MPORT_14_en = _T_162 & _GEN_15391;
  assign rf_MPORT_15_data = io_top_wb_bits_tc0_octet1_threadgroup4_matrix_d_data[63:0];
  assign rf_MPORT_15_addr = 8'he9;
  assign rf_MPORT_15_mask = 1'h1;
  assign rf_MPORT_15_en = _T_162 & _GEN_15391;
  assign rf_MPORT_16_data = io_top_wb_bits_tc1_octet0_threadgroup0_matrix_d_data[255:192];
  assign rf_MPORT_16_addr = 8'h84;
  assign rf_MPORT_16_mask = 1'h1;
  assign rf_MPORT_16_en = _T_162 & _GEN_15391;
  assign rf_MPORT_17_data = io_top_wb_bits_tc1_octet0_threadgroup0_matrix_d_data[191:128];
  assign rf_MPORT_17_addr = 8'h85;
  assign rf_MPORT_17_mask = 1'h1;
  assign rf_MPORT_17_en = _T_162 & _GEN_15391;
  assign rf_MPORT_18_data = io_top_wb_bits_tc1_octet0_threadgroup0_matrix_d_data[127:64];
  assign rf_MPORT_18_addr = 8'h8c;
  assign rf_MPORT_18_mask = 1'h1;
  assign rf_MPORT_18_en = _T_162 & _GEN_15391;
  assign rf_MPORT_19_data = io_top_wb_bits_tc1_octet0_threadgroup0_matrix_d_data[63:0];
  assign rf_MPORT_19_addr = 8'h8d;
  assign rf_MPORT_19_mask = 1'h1;
  assign rf_MPORT_19_en = _T_162 & _GEN_15391;
  assign rf_MPORT_20_data = io_top_wb_bits_tc1_octet0_threadgroup4_matrix_d_data[255:192];
  assign rf_MPORT_20_addr = 8'ha4;
  assign rf_MPORT_20_mask = 1'h1;
  assign rf_MPORT_20_en = _T_162 & _GEN_15391;
  assign rf_MPORT_21_data = io_top_wb_bits_tc1_octet0_threadgroup4_matrix_d_data[191:128];
  assign rf_MPORT_21_addr = 8'ha5;
  assign rf_MPORT_21_mask = 1'h1;
  assign rf_MPORT_21_en = _T_162 & _GEN_15391;
  assign rf_MPORT_22_data = io_top_wb_bits_tc1_octet0_threadgroup4_matrix_d_data[127:64];
  assign rf_MPORT_22_addr = 8'hac;
  assign rf_MPORT_22_mask = 1'h1;
  assign rf_MPORT_22_en = _T_162 & _GEN_15391;
  assign rf_MPORT_23_data = io_top_wb_bits_tc1_octet0_threadgroup4_matrix_d_data[63:0];
  assign rf_MPORT_23_addr = 8'had;
  assign rf_MPORT_23_mask = 1'h1;
  assign rf_MPORT_23_en = _T_162 & _GEN_15391;
  assign rf_MPORT_24_data = io_top_wb_bits_tc1_octet1_threadgroup0_matrix_d_data[255:192];
  assign rf_MPORT_24_addr = 8'hc4;
  assign rf_MPORT_24_mask = 1'h1;
  assign rf_MPORT_24_en = _T_162 & _GEN_15391;
  assign rf_MPORT_25_data = io_top_wb_bits_tc1_octet1_threadgroup0_matrix_d_data[191:128];
  assign rf_MPORT_25_addr = 8'hc5;
  assign rf_MPORT_25_mask = 1'h1;
  assign rf_MPORT_25_en = _T_162 & _GEN_15391;
  assign rf_MPORT_26_data = io_top_wb_bits_tc1_octet1_threadgroup0_matrix_d_data[127:64];
  assign rf_MPORT_26_addr = 8'hcc;
  assign rf_MPORT_26_mask = 1'h1;
  assign rf_MPORT_26_en = _T_162 & _GEN_15391;
  assign rf_MPORT_27_data = io_top_wb_bits_tc1_octet1_threadgroup0_matrix_d_data[63:0];
  assign rf_MPORT_27_addr = 8'hcd;
  assign rf_MPORT_27_mask = 1'h1;
  assign rf_MPORT_27_en = _T_162 & _GEN_15391;
  assign rf_MPORT_28_data = io_top_wb_bits_tc1_octet1_threadgroup4_matrix_d_data[255:192];
  assign rf_MPORT_28_addr = 8'he4;
  assign rf_MPORT_28_mask = 1'h1;
  assign rf_MPORT_28_en = _T_162 & _GEN_15391;
  assign rf_MPORT_29_data = io_top_wb_bits_tc1_octet1_threadgroup4_matrix_d_data[191:128];
  assign rf_MPORT_29_addr = 8'he5;
  assign rf_MPORT_29_mask = 1'h1;
  assign rf_MPORT_29_en = _T_162 & _GEN_15391;
  assign rf_MPORT_30_data = io_top_wb_bits_tc1_octet1_threadgroup4_matrix_d_data[127:64];
  assign rf_MPORT_30_addr = 8'hec;
  assign rf_MPORT_30_mask = 1'h1;
  assign rf_MPORT_30_en = _T_162 & _GEN_15391;
  assign rf_MPORT_31_data = io_top_wb_bits_tc1_octet1_threadgroup4_matrix_d_data[63:0];
  assign rf_MPORT_31_addr = 8'hed;
  assign rf_MPORT_31_mask = 1'h1;
  assign rf_MPORT_31_en = _T_162 & _GEN_15391;
  assign rf_MPORT_32_data = io_top_wb_bits_tc0_octet0_threadgroup0_matrix_d_data[255:192];
  assign rf_MPORT_32_addr = 8'h80;
  assign rf_MPORT_32_mask = 1'h1;
  assign rf_MPORT_32_en = _T_162 & _GEN_15458;
  assign rf_MPORT_33_data = io_top_wb_bits_tc0_octet0_threadgroup0_matrix_d_data[191:128];
  assign rf_MPORT_33_addr = 8'h84;
  assign rf_MPORT_33_mask = 1'h1;
  assign rf_MPORT_33_en = _T_162 & _GEN_15458;
  assign rf_MPORT_34_data = io_top_wb_bits_tc0_octet0_threadgroup0_matrix_d_data[127:64];
  assign rf_MPORT_34_addr = 8'h88;
  assign rf_MPORT_34_mask = 1'h1;
  assign rf_MPORT_34_en = _T_162 & _GEN_15458;
  assign rf_MPORT_35_data = io_top_wb_bits_tc0_octet0_threadgroup0_matrix_d_data[63:0];
  assign rf_MPORT_35_addr = 8'h8c;
  assign rf_MPORT_35_mask = 1'h1;
  assign rf_MPORT_35_en = _T_162 & _GEN_15458;
  assign rf_MPORT_36_data = io_top_wb_bits_tc0_octet0_threadgroup4_matrix_d_data[255:192];
  assign rf_MPORT_36_addr = 8'h90;
  assign rf_MPORT_36_mask = 1'h1;
  assign rf_MPORT_36_en = _T_162 & _GEN_15458;
  assign rf_MPORT_37_data = io_top_wb_bits_tc0_octet0_threadgroup4_matrix_d_data[191:128];
  assign rf_MPORT_37_addr = 8'h94;
  assign rf_MPORT_37_mask = 1'h1;
  assign rf_MPORT_37_en = _T_162 & _GEN_15458;
  assign rf_MPORT_38_data = io_top_wb_bits_tc0_octet0_threadgroup4_matrix_d_data[127:64];
  assign rf_MPORT_38_addr = 8'h98;
  assign rf_MPORT_38_mask = 1'h1;
  assign rf_MPORT_38_en = _T_162 & _GEN_15458;
  assign rf_MPORT_39_data = io_top_wb_bits_tc0_octet0_threadgroup4_matrix_d_data[63:0];
  assign rf_MPORT_39_addr = 8'h9c;
  assign rf_MPORT_39_mask = 1'h1;
  assign rf_MPORT_39_en = _T_162 & _GEN_15458;
  assign rf_MPORT_40_data = io_top_wb_bits_tc0_octet1_threadgroup0_matrix_d_data[255:192];
  assign rf_MPORT_40_addr = 8'ha0;
  assign rf_MPORT_40_mask = 1'h1;
  assign rf_MPORT_40_en = _T_162 & _GEN_15458;
  assign rf_MPORT_41_data = io_top_wb_bits_tc0_octet1_threadgroup0_matrix_d_data[191:128];
  assign rf_MPORT_41_addr = 8'ha4;
  assign rf_MPORT_41_mask = 1'h1;
  assign rf_MPORT_41_en = _T_162 & _GEN_15458;
  assign rf_MPORT_42_data = io_top_wb_bits_tc0_octet1_threadgroup0_matrix_d_data[127:64];
  assign rf_MPORT_42_addr = 8'ha8;
  assign rf_MPORT_42_mask = 1'h1;
  assign rf_MPORT_42_en = _T_162 & _GEN_15458;
  assign rf_MPORT_43_data = io_top_wb_bits_tc0_octet1_threadgroup0_matrix_d_data[63:0];
  assign rf_MPORT_43_addr = 8'hac;
  assign rf_MPORT_43_mask = 1'h1;
  assign rf_MPORT_43_en = _T_162 & _GEN_15458;
  assign rf_MPORT_44_data = io_top_wb_bits_tc0_octet1_threadgroup4_matrix_d_data[255:192];
  assign rf_MPORT_44_addr = 8'hb0;
  assign rf_MPORT_44_mask = 1'h1;
  assign rf_MPORT_44_en = _T_162 & _GEN_15458;
  assign rf_MPORT_45_data = io_top_wb_bits_tc0_octet1_threadgroup4_matrix_d_data[191:128];
  assign rf_MPORT_45_addr = 8'hb4;
  assign rf_MPORT_45_mask = 1'h1;
  assign rf_MPORT_45_en = _T_162 & _GEN_15458;
  assign rf_MPORT_46_data = io_top_wb_bits_tc0_octet1_threadgroup4_matrix_d_data[127:64];
  assign rf_MPORT_46_addr = 8'hb8;
  assign rf_MPORT_46_mask = 1'h1;
  assign rf_MPORT_46_en = _T_162 & _GEN_15458;
  assign rf_MPORT_47_data = io_top_wb_bits_tc0_octet1_threadgroup4_matrix_d_data[63:0];
  assign rf_MPORT_47_addr = 8'hbc;
  assign rf_MPORT_47_mask = 1'h1;
  assign rf_MPORT_47_en = _T_162 & _GEN_15458;
  assign rf_MPORT_48_data = io_top_wb_bits_tc1_octet0_threadgroup0_matrix_d_data[255:192];
  assign rf_MPORT_48_addr = 8'h82;
  assign rf_MPORT_48_mask = 1'h1;
  assign rf_MPORT_48_en = _T_162 & _GEN_15458;
  assign rf_MPORT_49_data = io_top_wb_bits_tc1_octet0_threadgroup0_matrix_d_data[191:128];
  assign rf_MPORT_49_addr = 8'h86;
  assign rf_MPORT_49_mask = 1'h1;
  assign rf_MPORT_49_en = _T_162 & _GEN_15458;
  assign rf_MPORT_50_data = io_top_wb_bits_tc1_octet0_threadgroup0_matrix_d_data[127:64];
  assign rf_MPORT_50_addr = 8'h8a;
  assign rf_MPORT_50_mask = 1'h1;
  assign rf_MPORT_50_en = _T_162 & _GEN_15458;
  assign rf_MPORT_51_data = io_top_wb_bits_tc1_octet0_threadgroup0_matrix_d_data[63:0];
  assign rf_MPORT_51_addr = 8'h8e;
  assign rf_MPORT_51_mask = 1'h1;
  assign rf_MPORT_51_en = _T_162 & _GEN_15458;
  assign rf_MPORT_52_data = io_top_wb_bits_tc1_octet0_threadgroup4_matrix_d_data[255:192];
  assign rf_MPORT_52_addr = 8'h92;
  assign rf_MPORT_52_mask = 1'h1;
  assign rf_MPORT_52_en = _T_162 & _GEN_15458;
  assign rf_MPORT_53_data = io_top_wb_bits_tc1_octet0_threadgroup4_matrix_d_data[191:128];
  assign rf_MPORT_53_addr = 8'h96;
  assign rf_MPORT_53_mask = 1'h1;
  assign rf_MPORT_53_en = _T_162 & _GEN_15458;
  assign rf_MPORT_54_data = io_top_wb_bits_tc1_octet0_threadgroup4_matrix_d_data[127:64];
  assign rf_MPORT_54_addr = 8'h9a;
  assign rf_MPORT_54_mask = 1'h1;
  assign rf_MPORT_54_en = _T_162 & _GEN_15458;
  assign rf_MPORT_55_data = io_top_wb_bits_tc1_octet0_threadgroup4_matrix_d_data[63:0];
  assign rf_MPORT_55_addr = 8'h9e;
  assign rf_MPORT_55_mask = 1'h1;
  assign rf_MPORT_55_en = _T_162 & _GEN_15458;
  assign rf_MPORT_56_data = io_top_wb_bits_tc1_octet1_threadgroup0_matrix_d_data[255:192];
  assign rf_MPORT_56_addr = 8'ha2;
  assign rf_MPORT_56_mask = 1'h1;
  assign rf_MPORT_56_en = _T_162 & _GEN_15458;
  assign rf_MPORT_57_data = io_top_wb_bits_tc1_octet1_threadgroup0_matrix_d_data[191:128];
  assign rf_MPORT_57_addr = 8'ha6;
  assign rf_MPORT_57_mask = 1'h1;
  assign rf_MPORT_57_en = _T_162 & _GEN_15458;
  assign rf_MPORT_58_data = io_top_wb_bits_tc1_octet1_threadgroup0_matrix_d_data[127:64];
  assign rf_MPORT_58_addr = 8'haa;
  assign rf_MPORT_58_mask = 1'h1;
  assign rf_MPORT_58_en = _T_162 & _GEN_15458;
  assign rf_MPORT_59_data = io_top_wb_bits_tc1_octet1_threadgroup0_matrix_d_data[63:0];
  assign rf_MPORT_59_addr = 8'hae;
  assign rf_MPORT_59_mask = 1'h1;
  assign rf_MPORT_59_en = _T_162 & _GEN_15458;
  assign rf_MPORT_60_data = io_top_wb_bits_tc1_octet1_threadgroup4_matrix_d_data[255:192];
  assign rf_MPORT_60_addr = 8'hb2;
  assign rf_MPORT_60_mask = 1'h1;
  assign rf_MPORT_60_en = _T_162 & _GEN_15458;
  assign rf_MPORT_61_data = io_top_wb_bits_tc1_octet1_threadgroup4_matrix_d_data[191:128];
  assign rf_MPORT_61_addr = 8'hb6;
  assign rf_MPORT_61_mask = 1'h1;
  assign rf_MPORT_61_en = _T_162 & _GEN_15458;
  assign rf_MPORT_62_data = io_top_wb_bits_tc1_octet1_threadgroup4_matrix_d_data[127:64];
  assign rf_MPORT_62_addr = 8'hba;
  assign rf_MPORT_62_mask = 1'h1;
  assign rf_MPORT_62_en = _T_162 & _GEN_15458;
  assign rf_MPORT_63_data = io_top_wb_bits_tc1_octet1_threadgroup4_matrix_d_data[63:0];
  assign rf_MPORT_63_addr = 8'hbe;
  assign rf_MPORT_63_mask = 1'h1;
  assign rf_MPORT_63_en = _T_162 & _GEN_15458;
  assign rf_MPORT_64_data = io_top_wb_bits_tc0_octet0_threadgroup0_matrix_d_data[255:192];
  assign rf_MPORT_64_addr = 8'h90;
  assign rf_MPORT_64_mask = 1'h1;
  assign rf_MPORT_64_en = _T_162 & _GEN_15525;
  assign rf_MPORT_65_data = io_top_wb_bits_tc0_octet0_threadgroup0_matrix_d_data[191:128];
  assign rf_MPORT_65_addr = 8'h91;
  assign rf_MPORT_65_mask = 1'h1;
  assign rf_MPORT_65_en = _T_162 & _GEN_15525;
  assign rf_MPORT_66_data = io_top_wb_bits_tc0_octet0_threadgroup0_matrix_d_data[127:64];
  assign rf_MPORT_66_addr = 8'h98;
  assign rf_MPORT_66_mask = 1'h1;
  assign rf_MPORT_66_en = _T_162 & _GEN_15525;
  assign rf_MPORT_67_data = io_top_wb_bits_tc0_octet0_threadgroup0_matrix_d_data[63:0];
  assign rf_MPORT_67_addr = 8'h99;
  assign rf_MPORT_67_mask = 1'h1;
  assign rf_MPORT_67_en = _T_162 & _GEN_15525;
  assign rf_MPORT_68_data = io_top_wb_bits_tc0_octet0_threadgroup4_matrix_d_data[255:192];
  assign rf_MPORT_68_addr = 8'hb0;
  assign rf_MPORT_68_mask = 1'h1;
  assign rf_MPORT_68_en = _T_162 & _GEN_15525;
  assign rf_MPORT_69_data = io_top_wb_bits_tc0_octet0_threadgroup4_matrix_d_data[191:128];
  assign rf_MPORT_69_addr = 8'hb1;
  assign rf_MPORT_69_mask = 1'h1;
  assign rf_MPORT_69_en = _T_162 & _GEN_15525;
  assign rf_MPORT_70_data = io_top_wb_bits_tc0_octet0_threadgroup4_matrix_d_data[127:64];
  assign rf_MPORT_70_addr = 8'hb8;
  assign rf_MPORT_70_mask = 1'h1;
  assign rf_MPORT_70_en = _T_162 & _GEN_15525;
  assign rf_MPORT_71_data = io_top_wb_bits_tc0_octet0_threadgroup4_matrix_d_data[63:0];
  assign rf_MPORT_71_addr = 8'hb9;
  assign rf_MPORT_71_mask = 1'h1;
  assign rf_MPORT_71_en = _T_162 & _GEN_15525;
  assign rf_MPORT_72_data = io_top_wb_bits_tc0_octet1_threadgroup0_matrix_d_data[255:192];
  assign rf_MPORT_72_addr = 8'hd0;
  assign rf_MPORT_72_mask = 1'h1;
  assign rf_MPORT_72_en = _T_162 & _GEN_15525;
  assign rf_MPORT_73_data = io_top_wb_bits_tc0_octet1_threadgroup0_matrix_d_data[191:128];
  assign rf_MPORT_73_addr = 8'hd1;
  assign rf_MPORT_73_mask = 1'h1;
  assign rf_MPORT_73_en = _T_162 & _GEN_15525;
  assign rf_MPORT_74_data = io_top_wb_bits_tc0_octet1_threadgroup0_matrix_d_data[127:64];
  assign rf_MPORT_74_addr = 8'hd8;
  assign rf_MPORT_74_mask = 1'h1;
  assign rf_MPORT_74_en = _T_162 & _GEN_15525;
  assign rf_MPORT_75_data = io_top_wb_bits_tc0_octet1_threadgroup0_matrix_d_data[63:0];
  assign rf_MPORT_75_addr = 8'hd9;
  assign rf_MPORT_75_mask = 1'h1;
  assign rf_MPORT_75_en = _T_162 & _GEN_15525;
  assign rf_MPORT_76_data = io_top_wb_bits_tc0_octet1_threadgroup4_matrix_d_data[255:192];
  assign rf_MPORT_76_addr = 8'hf0;
  assign rf_MPORT_76_mask = 1'h1;
  assign rf_MPORT_76_en = _T_162 & _GEN_15525;
  assign rf_MPORT_77_data = io_top_wb_bits_tc0_octet1_threadgroup4_matrix_d_data[191:128];
  assign rf_MPORT_77_addr = 8'hf1;
  assign rf_MPORT_77_mask = 1'h1;
  assign rf_MPORT_77_en = _T_162 & _GEN_15525;
  assign rf_MPORT_78_data = io_top_wb_bits_tc0_octet1_threadgroup4_matrix_d_data[127:64];
  assign rf_MPORT_78_addr = 8'hf8;
  assign rf_MPORT_78_mask = 1'h1;
  assign rf_MPORT_78_en = _T_162 & _GEN_15525;
  assign rf_MPORT_79_data = io_top_wb_bits_tc0_octet1_threadgroup4_matrix_d_data[63:0];
  assign rf_MPORT_79_addr = 8'hf9;
  assign rf_MPORT_79_mask = 1'h1;
  assign rf_MPORT_79_en = _T_162 & _GEN_15525;
  assign rf_MPORT_80_data = io_top_wb_bits_tc1_octet0_threadgroup0_matrix_d_data[255:192];
  assign rf_MPORT_80_addr = 8'h94;
  assign rf_MPORT_80_mask = 1'h1;
  assign rf_MPORT_80_en = _T_162 & _GEN_15525;
  assign rf_MPORT_81_data = io_top_wb_bits_tc1_octet0_threadgroup0_matrix_d_data[191:128];
  assign rf_MPORT_81_addr = 8'h95;
  assign rf_MPORT_81_mask = 1'h1;
  assign rf_MPORT_81_en = _T_162 & _GEN_15525;
  assign rf_MPORT_82_data = io_top_wb_bits_tc1_octet0_threadgroup0_matrix_d_data[127:64];
  assign rf_MPORT_82_addr = 8'h9c;
  assign rf_MPORT_82_mask = 1'h1;
  assign rf_MPORT_82_en = _T_162 & _GEN_15525;
  assign rf_MPORT_83_data = io_top_wb_bits_tc1_octet0_threadgroup0_matrix_d_data[63:0];
  assign rf_MPORT_83_addr = 8'h9d;
  assign rf_MPORT_83_mask = 1'h1;
  assign rf_MPORT_83_en = _T_162 & _GEN_15525;
  assign rf_MPORT_84_data = io_top_wb_bits_tc1_octet0_threadgroup4_matrix_d_data[255:192];
  assign rf_MPORT_84_addr = 8'hb4;
  assign rf_MPORT_84_mask = 1'h1;
  assign rf_MPORT_84_en = _T_162 & _GEN_15525;
  assign rf_MPORT_85_data = io_top_wb_bits_tc1_octet0_threadgroup4_matrix_d_data[191:128];
  assign rf_MPORT_85_addr = 8'hb5;
  assign rf_MPORT_85_mask = 1'h1;
  assign rf_MPORT_85_en = _T_162 & _GEN_15525;
  assign rf_MPORT_86_data = io_top_wb_bits_tc1_octet0_threadgroup4_matrix_d_data[127:64];
  assign rf_MPORT_86_addr = 8'hbc;
  assign rf_MPORT_86_mask = 1'h1;
  assign rf_MPORT_86_en = _T_162 & _GEN_15525;
  assign rf_MPORT_87_data = io_top_wb_bits_tc1_octet0_threadgroup4_matrix_d_data[63:0];
  assign rf_MPORT_87_addr = 8'hbd;
  assign rf_MPORT_87_mask = 1'h1;
  assign rf_MPORT_87_en = _T_162 & _GEN_15525;
  assign rf_MPORT_88_data = io_top_wb_bits_tc1_octet1_threadgroup0_matrix_d_data[255:192];
  assign rf_MPORT_88_addr = 8'hd4;
  assign rf_MPORT_88_mask = 1'h1;
  assign rf_MPORT_88_en = _T_162 & _GEN_15525;
  assign rf_MPORT_89_data = io_top_wb_bits_tc1_octet1_threadgroup0_matrix_d_data[191:128];
  assign rf_MPORT_89_addr = 8'hd5;
  assign rf_MPORT_89_mask = 1'h1;
  assign rf_MPORT_89_en = _T_162 & _GEN_15525;
  assign rf_MPORT_90_data = io_top_wb_bits_tc1_octet1_threadgroup0_matrix_d_data[127:64];
  assign rf_MPORT_90_addr = 8'hdc;
  assign rf_MPORT_90_mask = 1'h1;
  assign rf_MPORT_90_en = _T_162 & _GEN_15525;
  assign rf_MPORT_91_data = io_top_wb_bits_tc1_octet1_threadgroup0_matrix_d_data[63:0];
  assign rf_MPORT_91_addr = 8'hdd;
  assign rf_MPORT_91_mask = 1'h1;
  assign rf_MPORT_91_en = _T_162 & _GEN_15525;
  assign rf_MPORT_92_data = io_top_wb_bits_tc1_octet1_threadgroup4_matrix_d_data[255:192];
  assign rf_MPORT_92_addr = 8'hf4;
  assign rf_MPORT_92_mask = 1'h1;
  assign rf_MPORT_92_en = _T_162 & _GEN_15525;
  assign rf_MPORT_93_data = io_top_wb_bits_tc1_octet1_threadgroup4_matrix_d_data[191:128];
  assign rf_MPORT_93_addr = 8'hf5;
  assign rf_MPORT_93_mask = 1'h1;
  assign rf_MPORT_93_en = _T_162 & _GEN_15525;
  assign rf_MPORT_94_data = io_top_wb_bits_tc1_octet1_threadgroup4_matrix_d_data[127:64];
  assign rf_MPORT_94_addr = 8'hfc;
  assign rf_MPORT_94_mask = 1'h1;
  assign rf_MPORT_94_en = _T_162 & _GEN_15525;
  assign rf_MPORT_95_data = io_top_wb_bits_tc1_octet1_threadgroup4_matrix_d_data[63:0];
  assign rf_MPORT_95_addr = 8'hfd;
  assign rf_MPORT_95_mask = 1'h1;
  assign rf_MPORT_95_en = _T_162 & _GEN_15525;
  assign rf_MPORT_96_data = io_top_wb_bits_tc0_octet0_threadgroup0_matrix_d_data[255:192];
  assign rf_MPORT_96_addr = 8'h81;
  assign rf_MPORT_96_mask = 1'h1;
  assign rf_MPORT_96_en = _T_162 & _GEN_15592;
  assign rf_MPORT_97_data = io_top_wb_bits_tc0_octet0_threadgroup0_matrix_d_data[191:128];
  assign rf_MPORT_97_addr = 8'h85;
  assign rf_MPORT_97_mask = 1'h1;
  assign rf_MPORT_97_en = _T_162 & _GEN_15592;
  assign rf_MPORT_98_data = io_top_wb_bits_tc0_octet0_threadgroup0_matrix_d_data[127:64];
  assign rf_MPORT_98_addr = 8'h89;
  assign rf_MPORT_98_mask = 1'h1;
  assign rf_MPORT_98_en = _T_162 & _GEN_15592;
  assign rf_MPORT_99_data = io_top_wb_bits_tc0_octet0_threadgroup0_matrix_d_data[63:0];
  assign rf_MPORT_99_addr = 8'h8d;
  assign rf_MPORT_99_mask = 1'h1;
  assign rf_MPORT_99_en = _T_162 & _GEN_15592;
  assign rf_MPORT_100_data = io_top_wb_bits_tc0_octet0_threadgroup4_matrix_d_data[255:192];
  assign rf_MPORT_100_addr = 8'h91;
  assign rf_MPORT_100_mask = 1'h1;
  assign rf_MPORT_100_en = _T_162 & _GEN_15592;
  assign rf_MPORT_101_data = io_top_wb_bits_tc0_octet0_threadgroup4_matrix_d_data[191:128];
  assign rf_MPORT_101_addr = 8'h95;
  assign rf_MPORT_101_mask = 1'h1;
  assign rf_MPORT_101_en = _T_162 & _GEN_15592;
  assign rf_MPORT_102_data = io_top_wb_bits_tc0_octet0_threadgroup4_matrix_d_data[127:64];
  assign rf_MPORT_102_addr = 8'h99;
  assign rf_MPORT_102_mask = 1'h1;
  assign rf_MPORT_102_en = _T_162 & _GEN_15592;
  assign rf_MPORT_103_data = io_top_wb_bits_tc0_octet0_threadgroup4_matrix_d_data[63:0];
  assign rf_MPORT_103_addr = 8'h9d;
  assign rf_MPORT_103_mask = 1'h1;
  assign rf_MPORT_103_en = _T_162 & _GEN_15592;
  assign rf_MPORT_104_data = io_top_wb_bits_tc0_octet1_threadgroup0_matrix_d_data[255:192];
  assign rf_MPORT_104_addr = 8'ha1;
  assign rf_MPORT_104_mask = 1'h1;
  assign rf_MPORT_104_en = _T_162 & _GEN_15592;
  assign rf_MPORT_105_data = io_top_wb_bits_tc0_octet1_threadgroup0_matrix_d_data[191:128];
  assign rf_MPORT_105_addr = 8'ha5;
  assign rf_MPORT_105_mask = 1'h1;
  assign rf_MPORT_105_en = _T_162 & _GEN_15592;
  assign rf_MPORT_106_data = io_top_wb_bits_tc0_octet1_threadgroup0_matrix_d_data[127:64];
  assign rf_MPORT_106_addr = 8'ha9;
  assign rf_MPORT_106_mask = 1'h1;
  assign rf_MPORT_106_en = _T_162 & _GEN_15592;
  assign rf_MPORT_107_data = io_top_wb_bits_tc0_octet1_threadgroup0_matrix_d_data[63:0];
  assign rf_MPORT_107_addr = 8'had;
  assign rf_MPORT_107_mask = 1'h1;
  assign rf_MPORT_107_en = _T_162 & _GEN_15592;
  assign rf_MPORT_108_data = io_top_wb_bits_tc0_octet1_threadgroup4_matrix_d_data[255:192];
  assign rf_MPORT_108_addr = 8'hb1;
  assign rf_MPORT_108_mask = 1'h1;
  assign rf_MPORT_108_en = _T_162 & _GEN_15592;
  assign rf_MPORT_109_data = io_top_wb_bits_tc0_octet1_threadgroup4_matrix_d_data[191:128];
  assign rf_MPORT_109_addr = 8'hb5;
  assign rf_MPORT_109_mask = 1'h1;
  assign rf_MPORT_109_en = _T_162 & _GEN_15592;
  assign rf_MPORT_110_data = io_top_wb_bits_tc0_octet1_threadgroup4_matrix_d_data[127:64];
  assign rf_MPORT_110_addr = 8'hb9;
  assign rf_MPORT_110_mask = 1'h1;
  assign rf_MPORT_110_en = _T_162 & _GEN_15592;
  assign rf_MPORT_111_data = io_top_wb_bits_tc0_octet1_threadgroup4_matrix_d_data[63:0];
  assign rf_MPORT_111_addr = 8'hbd;
  assign rf_MPORT_111_mask = 1'h1;
  assign rf_MPORT_111_en = _T_162 & _GEN_15592;
  assign rf_MPORT_112_data = io_top_wb_bits_tc1_octet0_threadgroup0_matrix_d_data[255:192];
  assign rf_MPORT_112_addr = 8'h83;
  assign rf_MPORT_112_mask = 1'h1;
  assign rf_MPORT_112_en = _T_162 & _GEN_15592;
  assign rf_MPORT_113_data = io_top_wb_bits_tc1_octet0_threadgroup0_matrix_d_data[191:128];
  assign rf_MPORT_113_addr = 8'h87;
  assign rf_MPORT_113_mask = 1'h1;
  assign rf_MPORT_113_en = _T_162 & _GEN_15592;
  assign rf_MPORT_114_data = io_top_wb_bits_tc1_octet0_threadgroup0_matrix_d_data[127:64];
  assign rf_MPORT_114_addr = 8'h8b;
  assign rf_MPORT_114_mask = 1'h1;
  assign rf_MPORT_114_en = _T_162 & _GEN_15592;
  assign rf_MPORT_115_data = io_top_wb_bits_tc1_octet0_threadgroup0_matrix_d_data[63:0];
  assign rf_MPORT_115_addr = 8'h8f;
  assign rf_MPORT_115_mask = 1'h1;
  assign rf_MPORT_115_en = _T_162 & _GEN_15592;
  assign rf_MPORT_116_data = io_top_wb_bits_tc1_octet0_threadgroup4_matrix_d_data[255:192];
  assign rf_MPORT_116_addr = 8'h93;
  assign rf_MPORT_116_mask = 1'h1;
  assign rf_MPORT_116_en = _T_162 & _GEN_15592;
  assign rf_MPORT_117_data = io_top_wb_bits_tc1_octet0_threadgroup4_matrix_d_data[191:128];
  assign rf_MPORT_117_addr = 8'h97;
  assign rf_MPORT_117_mask = 1'h1;
  assign rf_MPORT_117_en = _T_162 & _GEN_15592;
  assign rf_MPORT_118_data = io_top_wb_bits_tc1_octet0_threadgroup4_matrix_d_data[127:64];
  assign rf_MPORT_118_addr = 8'h9b;
  assign rf_MPORT_118_mask = 1'h1;
  assign rf_MPORT_118_en = _T_162 & _GEN_15592;
  assign rf_MPORT_119_data = io_top_wb_bits_tc1_octet0_threadgroup4_matrix_d_data[63:0];
  assign rf_MPORT_119_addr = 8'h9f;
  assign rf_MPORT_119_mask = 1'h1;
  assign rf_MPORT_119_en = _T_162 & _GEN_15592;
  assign rf_MPORT_120_data = io_top_wb_bits_tc1_octet1_threadgroup0_matrix_d_data[255:192];
  assign rf_MPORT_120_addr = 8'ha3;
  assign rf_MPORT_120_mask = 1'h1;
  assign rf_MPORT_120_en = _T_162 & _GEN_15592;
  assign rf_MPORT_121_data = io_top_wb_bits_tc1_octet1_threadgroup0_matrix_d_data[191:128];
  assign rf_MPORT_121_addr = 8'ha7;
  assign rf_MPORT_121_mask = 1'h1;
  assign rf_MPORT_121_en = _T_162 & _GEN_15592;
  assign rf_MPORT_122_data = io_top_wb_bits_tc1_octet1_threadgroup0_matrix_d_data[127:64];
  assign rf_MPORT_122_addr = 8'hab;
  assign rf_MPORT_122_mask = 1'h1;
  assign rf_MPORT_122_en = _T_162 & _GEN_15592;
  assign rf_MPORT_123_data = io_top_wb_bits_tc1_octet1_threadgroup0_matrix_d_data[63:0];
  assign rf_MPORT_123_addr = 8'haf;
  assign rf_MPORT_123_mask = 1'h1;
  assign rf_MPORT_123_en = _T_162 & _GEN_15592;
  assign rf_MPORT_124_data = io_top_wb_bits_tc1_octet1_threadgroup4_matrix_d_data[255:192];
  assign rf_MPORT_124_addr = 8'hb3;
  assign rf_MPORT_124_mask = 1'h1;
  assign rf_MPORT_124_en = _T_162 & _GEN_15592;
  assign rf_MPORT_125_data = io_top_wb_bits_tc1_octet1_threadgroup4_matrix_d_data[191:128];
  assign rf_MPORT_125_addr = 8'hb7;
  assign rf_MPORT_125_mask = 1'h1;
  assign rf_MPORT_125_en = _T_162 & _GEN_15592;
  assign rf_MPORT_126_data = io_top_wb_bits_tc1_octet1_threadgroup4_matrix_d_data[127:64];
  assign rf_MPORT_126_addr = 8'hbb;
  assign rf_MPORT_126_mask = 1'h1;
  assign rf_MPORT_126_en = _T_162 & _GEN_15592;
  assign rf_MPORT_127_data = io_top_wb_bits_tc1_octet1_threadgroup4_matrix_d_data[63:0];
  assign rf_MPORT_127_addr = 8'hbf;
  assign rf_MPORT_127_mask = 1'h1;
  assign rf_MPORT_127_en = _T_162 & _GEN_15592;
  assign rf_MPORT_128_data = io_top_wb_bits_tc0_octet0_threadgroup0_matrix_d_data[255:192];
  assign rf_MPORT_128_addr = 8'h82;
  assign rf_MPORT_128_mask = 1'h1;
  assign rf_MPORT_128_en = _T_162 & _GEN_15659;
  assign rf_MPORT_129_data = io_top_wb_bits_tc0_octet0_threadgroup0_matrix_d_data[191:128];
  assign rf_MPORT_129_addr = 8'h83;
  assign rf_MPORT_129_mask = 1'h1;
  assign rf_MPORT_129_en = _T_162 & _GEN_15659;
  assign rf_MPORT_130_data = io_top_wb_bits_tc0_octet0_threadgroup0_matrix_d_data[127:64];
  assign rf_MPORT_130_addr = 8'h8a;
  assign rf_MPORT_130_mask = 1'h1;
  assign rf_MPORT_130_en = _T_162 & _GEN_15659;
  assign rf_MPORT_131_data = io_top_wb_bits_tc0_octet0_threadgroup0_matrix_d_data[63:0];
  assign rf_MPORT_131_addr = 8'h8b;
  assign rf_MPORT_131_mask = 1'h1;
  assign rf_MPORT_131_en = _T_162 & _GEN_15659;
  assign rf_MPORT_132_data = io_top_wb_bits_tc0_octet0_threadgroup4_matrix_d_data[255:192];
  assign rf_MPORT_132_addr = 8'ha2;
  assign rf_MPORT_132_mask = 1'h1;
  assign rf_MPORT_132_en = _T_162 & _GEN_15659;
  assign rf_MPORT_133_data = io_top_wb_bits_tc0_octet0_threadgroup4_matrix_d_data[191:128];
  assign rf_MPORT_133_addr = 8'ha3;
  assign rf_MPORT_133_mask = 1'h1;
  assign rf_MPORT_133_en = _T_162 & _GEN_15659;
  assign rf_MPORT_134_data = io_top_wb_bits_tc0_octet0_threadgroup4_matrix_d_data[127:64];
  assign rf_MPORT_134_addr = 8'haa;
  assign rf_MPORT_134_mask = 1'h1;
  assign rf_MPORT_134_en = _T_162 & _GEN_15659;
  assign rf_MPORT_135_data = io_top_wb_bits_tc0_octet0_threadgroup4_matrix_d_data[63:0];
  assign rf_MPORT_135_addr = 8'hab;
  assign rf_MPORT_135_mask = 1'h1;
  assign rf_MPORT_135_en = _T_162 & _GEN_15659;
  assign rf_MPORT_136_data = io_top_wb_bits_tc0_octet1_threadgroup0_matrix_d_data[255:192];
  assign rf_MPORT_136_addr = 8'hc2;
  assign rf_MPORT_136_mask = 1'h1;
  assign rf_MPORT_136_en = _T_162 & _GEN_15659;
  assign rf_MPORT_137_data = io_top_wb_bits_tc0_octet1_threadgroup0_matrix_d_data[191:128];
  assign rf_MPORT_137_addr = 8'hc3;
  assign rf_MPORT_137_mask = 1'h1;
  assign rf_MPORT_137_en = _T_162 & _GEN_15659;
  assign rf_MPORT_138_data = io_top_wb_bits_tc0_octet1_threadgroup0_matrix_d_data[127:64];
  assign rf_MPORT_138_addr = 8'hca;
  assign rf_MPORT_138_mask = 1'h1;
  assign rf_MPORT_138_en = _T_162 & _GEN_15659;
  assign rf_MPORT_139_data = io_top_wb_bits_tc0_octet1_threadgroup0_matrix_d_data[63:0];
  assign rf_MPORT_139_addr = 8'hcb;
  assign rf_MPORT_139_mask = 1'h1;
  assign rf_MPORT_139_en = _T_162 & _GEN_15659;
  assign rf_MPORT_140_data = io_top_wb_bits_tc0_octet1_threadgroup4_matrix_d_data[255:192];
  assign rf_MPORT_140_addr = 8'he2;
  assign rf_MPORT_140_mask = 1'h1;
  assign rf_MPORT_140_en = _T_162 & _GEN_15659;
  assign rf_MPORT_141_data = io_top_wb_bits_tc0_octet1_threadgroup4_matrix_d_data[191:128];
  assign rf_MPORT_141_addr = 8'he3;
  assign rf_MPORT_141_mask = 1'h1;
  assign rf_MPORT_141_en = _T_162 & _GEN_15659;
  assign rf_MPORT_142_data = io_top_wb_bits_tc0_octet1_threadgroup4_matrix_d_data[127:64];
  assign rf_MPORT_142_addr = 8'hea;
  assign rf_MPORT_142_mask = 1'h1;
  assign rf_MPORT_142_en = _T_162 & _GEN_15659;
  assign rf_MPORT_143_data = io_top_wb_bits_tc0_octet1_threadgroup4_matrix_d_data[63:0];
  assign rf_MPORT_143_addr = 8'heb;
  assign rf_MPORT_143_mask = 1'h1;
  assign rf_MPORT_143_en = _T_162 & _GEN_15659;
  assign rf_MPORT_144_data = io_top_wb_bits_tc1_octet0_threadgroup0_matrix_d_data[255:192];
  assign rf_MPORT_144_addr = 8'h86;
  assign rf_MPORT_144_mask = 1'h1;
  assign rf_MPORT_144_en = _T_162 & _GEN_15659;
  assign rf_MPORT_145_data = io_top_wb_bits_tc1_octet0_threadgroup0_matrix_d_data[191:128];
  assign rf_MPORT_145_addr = 8'h87;
  assign rf_MPORT_145_mask = 1'h1;
  assign rf_MPORT_145_en = _T_162 & _GEN_15659;
  assign rf_MPORT_146_data = io_top_wb_bits_tc1_octet0_threadgroup0_matrix_d_data[127:64];
  assign rf_MPORT_146_addr = 8'h8e;
  assign rf_MPORT_146_mask = 1'h1;
  assign rf_MPORT_146_en = _T_162 & _GEN_15659;
  assign rf_MPORT_147_data = io_top_wb_bits_tc1_octet0_threadgroup0_matrix_d_data[63:0];
  assign rf_MPORT_147_addr = 8'h8f;
  assign rf_MPORT_147_mask = 1'h1;
  assign rf_MPORT_147_en = _T_162 & _GEN_15659;
  assign rf_MPORT_148_data = io_top_wb_bits_tc1_octet0_threadgroup4_matrix_d_data[255:192];
  assign rf_MPORT_148_addr = 8'ha6;
  assign rf_MPORT_148_mask = 1'h1;
  assign rf_MPORT_148_en = _T_162 & _GEN_15659;
  assign rf_MPORT_149_data = io_top_wb_bits_tc1_octet0_threadgroup4_matrix_d_data[191:128];
  assign rf_MPORT_149_addr = 8'ha7;
  assign rf_MPORT_149_mask = 1'h1;
  assign rf_MPORT_149_en = _T_162 & _GEN_15659;
  assign rf_MPORT_150_data = io_top_wb_bits_tc1_octet0_threadgroup4_matrix_d_data[127:64];
  assign rf_MPORT_150_addr = 8'hae;
  assign rf_MPORT_150_mask = 1'h1;
  assign rf_MPORT_150_en = _T_162 & _GEN_15659;
  assign rf_MPORT_151_data = io_top_wb_bits_tc1_octet0_threadgroup4_matrix_d_data[63:0];
  assign rf_MPORT_151_addr = 8'haf;
  assign rf_MPORT_151_mask = 1'h1;
  assign rf_MPORT_151_en = _T_162 & _GEN_15659;
  assign rf_MPORT_152_data = io_top_wb_bits_tc1_octet1_threadgroup0_matrix_d_data[255:192];
  assign rf_MPORT_152_addr = 8'hc6;
  assign rf_MPORT_152_mask = 1'h1;
  assign rf_MPORT_152_en = _T_162 & _GEN_15659;
  assign rf_MPORT_153_data = io_top_wb_bits_tc1_octet1_threadgroup0_matrix_d_data[191:128];
  assign rf_MPORT_153_addr = 8'hc7;
  assign rf_MPORT_153_mask = 1'h1;
  assign rf_MPORT_153_en = _T_162 & _GEN_15659;
  assign rf_MPORT_154_data = io_top_wb_bits_tc1_octet1_threadgroup0_matrix_d_data[127:64];
  assign rf_MPORT_154_addr = 8'hce;
  assign rf_MPORT_154_mask = 1'h1;
  assign rf_MPORT_154_en = _T_162 & _GEN_15659;
  assign rf_MPORT_155_data = io_top_wb_bits_tc1_octet1_threadgroup0_matrix_d_data[63:0];
  assign rf_MPORT_155_addr = 8'hcf;
  assign rf_MPORT_155_mask = 1'h1;
  assign rf_MPORT_155_en = _T_162 & _GEN_15659;
  assign rf_MPORT_156_data = io_top_wb_bits_tc1_octet1_threadgroup4_matrix_d_data[255:192];
  assign rf_MPORT_156_addr = 8'he6;
  assign rf_MPORT_156_mask = 1'h1;
  assign rf_MPORT_156_en = _T_162 & _GEN_15659;
  assign rf_MPORT_157_data = io_top_wb_bits_tc1_octet1_threadgroup4_matrix_d_data[191:128];
  assign rf_MPORT_157_addr = 8'he7;
  assign rf_MPORT_157_mask = 1'h1;
  assign rf_MPORT_157_en = _T_162 & _GEN_15659;
  assign rf_MPORT_158_data = io_top_wb_bits_tc1_octet1_threadgroup4_matrix_d_data[127:64];
  assign rf_MPORT_158_addr = 8'hee;
  assign rf_MPORT_158_mask = 1'h1;
  assign rf_MPORT_158_en = _T_162 & _GEN_15659;
  assign rf_MPORT_159_data = io_top_wb_bits_tc1_octet1_threadgroup4_matrix_d_data[63:0];
  assign rf_MPORT_159_addr = 8'hef;
  assign rf_MPORT_159_mask = 1'h1;
  assign rf_MPORT_159_en = _T_162 & _GEN_15659;
  assign rf_MPORT_160_data = io_top_wb_bits_tc0_octet0_threadgroup0_matrix_d_data[255:192];
  assign rf_MPORT_160_addr = 8'h92;
  assign rf_MPORT_160_mask = 1'h1;
  assign rf_MPORT_160_en = _T_162 & _GEN_15726;
  assign rf_MPORT_161_data = io_top_wb_bits_tc0_octet0_threadgroup0_matrix_d_data[191:128];
  assign rf_MPORT_161_addr = 8'h93;
  assign rf_MPORT_161_mask = 1'h1;
  assign rf_MPORT_161_en = _T_162 & _GEN_15726;
  assign rf_MPORT_162_data = io_top_wb_bits_tc0_octet0_threadgroup0_matrix_d_data[127:64];
  assign rf_MPORT_162_addr = 8'h9a;
  assign rf_MPORT_162_mask = 1'h1;
  assign rf_MPORT_162_en = _T_162 & _GEN_15726;
  assign rf_MPORT_163_data = io_top_wb_bits_tc0_octet0_threadgroup0_matrix_d_data[63:0];
  assign rf_MPORT_163_addr = 8'h9b;
  assign rf_MPORT_163_mask = 1'h1;
  assign rf_MPORT_163_en = _T_162 & _GEN_15726;
  assign rf_MPORT_164_data = io_top_wb_bits_tc0_octet0_threadgroup4_matrix_d_data[255:192];
  assign rf_MPORT_164_addr = 8'hb2;
  assign rf_MPORT_164_mask = 1'h1;
  assign rf_MPORT_164_en = _T_162 & _GEN_15726;
  assign rf_MPORT_165_data = io_top_wb_bits_tc0_octet0_threadgroup4_matrix_d_data[191:128];
  assign rf_MPORT_165_addr = 8'hb3;
  assign rf_MPORT_165_mask = 1'h1;
  assign rf_MPORT_165_en = _T_162 & _GEN_15726;
  assign rf_MPORT_166_data = io_top_wb_bits_tc0_octet0_threadgroup4_matrix_d_data[127:64];
  assign rf_MPORT_166_addr = 8'hba;
  assign rf_MPORT_166_mask = 1'h1;
  assign rf_MPORT_166_en = _T_162 & _GEN_15726;
  assign rf_MPORT_167_data = io_top_wb_bits_tc0_octet0_threadgroup4_matrix_d_data[63:0];
  assign rf_MPORT_167_addr = 8'hbb;
  assign rf_MPORT_167_mask = 1'h1;
  assign rf_MPORT_167_en = _T_162 & _GEN_15726;
  assign rf_MPORT_168_data = io_top_wb_bits_tc0_octet1_threadgroup0_matrix_d_data[255:192];
  assign rf_MPORT_168_addr = 8'hd2;
  assign rf_MPORT_168_mask = 1'h1;
  assign rf_MPORT_168_en = _T_162 & _GEN_15726;
  assign rf_MPORT_169_data = io_top_wb_bits_tc0_octet1_threadgroup0_matrix_d_data[191:128];
  assign rf_MPORT_169_addr = 8'hd3;
  assign rf_MPORT_169_mask = 1'h1;
  assign rf_MPORT_169_en = _T_162 & _GEN_15726;
  assign rf_MPORT_170_data = io_top_wb_bits_tc0_octet1_threadgroup0_matrix_d_data[127:64];
  assign rf_MPORT_170_addr = 8'hda;
  assign rf_MPORT_170_mask = 1'h1;
  assign rf_MPORT_170_en = _T_162 & _GEN_15726;
  assign rf_MPORT_171_data = io_top_wb_bits_tc0_octet1_threadgroup0_matrix_d_data[63:0];
  assign rf_MPORT_171_addr = 8'hdb;
  assign rf_MPORT_171_mask = 1'h1;
  assign rf_MPORT_171_en = _T_162 & _GEN_15726;
  assign rf_MPORT_172_data = io_top_wb_bits_tc0_octet1_threadgroup4_matrix_d_data[255:192];
  assign rf_MPORT_172_addr = 8'hf2;
  assign rf_MPORT_172_mask = 1'h1;
  assign rf_MPORT_172_en = _T_162 & _GEN_15726;
  assign rf_MPORT_173_data = io_top_wb_bits_tc0_octet1_threadgroup4_matrix_d_data[191:128];
  assign rf_MPORT_173_addr = 8'hf3;
  assign rf_MPORT_173_mask = 1'h1;
  assign rf_MPORT_173_en = _T_162 & _GEN_15726;
  assign rf_MPORT_174_data = io_top_wb_bits_tc0_octet1_threadgroup4_matrix_d_data[127:64];
  assign rf_MPORT_174_addr = 8'hfa;
  assign rf_MPORT_174_mask = 1'h1;
  assign rf_MPORT_174_en = _T_162 & _GEN_15726;
  assign rf_MPORT_175_data = io_top_wb_bits_tc0_octet1_threadgroup4_matrix_d_data[63:0];
  assign rf_MPORT_175_addr = 8'hfb;
  assign rf_MPORT_175_mask = 1'h1;
  assign rf_MPORT_175_en = _T_162 & _GEN_15726;
  assign rf_MPORT_176_data = io_top_wb_bits_tc1_octet0_threadgroup0_matrix_d_data[255:192];
  assign rf_MPORT_176_addr = 8'h96;
  assign rf_MPORT_176_mask = 1'h1;
  assign rf_MPORT_176_en = _T_162 & _GEN_15726;
  assign rf_MPORT_177_data = io_top_wb_bits_tc1_octet0_threadgroup0_matrix_d_data[191:128];
  assign rf_MPORT_177_addr = 8'h97;
  assign rf_MPORT_177_mask = 1'h1;
  assign rf_MPORT_177_en = _T_162 & _GEN_15726;
  assign rf_MPORT_178_data = io_top_wb_bits_tc1_octet0_threadgroup0_matrix_d_data[127:64];
  assign rf_MPORT_178_addr = 8'h9e;
  assign rf_MPORT_178_mask = 1'h1;
  assign rf_MPORT_178_en = _T_162 & _GEN_15726;
  assign rf_MPORT_179_data = io_top_wb_bits_tc1_octet0_threadgroup0_matrix_d_data[63:0];
  assign rf_MPORT_179_addr = 8'h9f;
  assign rf_MPORT_179_mask = 1'h1;
  assign rf_MPORT_179_en = _T_162 & _GEN_15726;
  assign rf_MPORT_180_data = io_top_wb_bits_tc1_octet0_threadgroup4_matrix_d_data[255:192];
  assign rf_MPORT_180_addr = 8'hb6;
  assign rf_MPORT_180_mask = 1'h1;
  assign rf_MPORT_180_en = _T_162 & _GEN_15726;
  assign rf_MPORT_181_data = io_top_wb_bits_tc1_octet0_threadgroup4_matrix_d_data[191:128];
  assign rf_MPORT_181_addr = 8'hb7;
  assign rf_MPORT_181_mask = 1'h1;
  assign rf_MPORT_181_en = _T_162 & _GEN_15726;
  assign rf_MPORT_182_data = io_top_wb_bits_tc1_octet0_threadgroup4_matrix_d_data[127:64];
  assign rf_MPORT_182_addr = 8'hbe;
  assign rf_MPORT_182_mask = 1'h1;
  assign rf_MPORT_182_en = _T_162 & _GEN_15726;
  assign rf_MPORT_183_data = io_top_wb_bits_tc1_octet0_threadgroup4_matrix_d_data[63:0];
  assign rf_MPORT_183_addr = 8'hbf;
  assign rf_MPORT_183_mask = 1'h1;
  assign rf_MPORT_183_en = _T_162 & _GEN_15726;
  assign rf_MPORT_184_data = io_top_wb_bits_tc1_octet1_threadgroup0_matrix_d_data[255:192];
  assign rf_MPORT_184_addr = 8'hd6;
  assign rf_MPORT_184_mask = 1'h1;
  assign rf_MPORT_184_en = _T_162 & _GEN_15726;
  assign rf_MPORT_185_data = io_top_wb_bits_tc1_octet1_threadgroup0_matrix_d_data[191:128];
  assign rf_MPORT_185_addr = 8'hd7;
  assign rf_MPORT_185_mask = 1'h1;
  assign rf_MPORT_185_en = _T_162 & _GEN_15726;
  assign rf_MPORT_186_data = io_top_wb_bits_tc1_octet1_threadgroup0_matrix_d_data[127:64];
  assign rf_MPORT_186_addr = 8'hde;
  assign rf_MPORT_186_mask = 1'h1;
  assign rf_MPORT_186_en = _T_162 & _GEN_15726;
  assign rf_MPORT_187_data = io_top_wb_bits_tc1_octet1_threadgroup0_matrix_d_data[63:0];
  assign rf_MPORT_187_addr = 8'hdf;
  assign rf_MPORT_187_mask = 1'h1;
  assign rf_MPORT_187_en = _T_162 & _GEN_15726;
  assign rf_MPORT_188_data = io_top_wb_bits_tc1_octet1_threadgroup4_matrix_d_data[255:192];
  assign rf_MPORT_188_addr = 8'hf6;
  assign rf_MPORT_188_mask = 1'h1;
  assign rf_MPORT_188_en = _T_162 & _GEN_15726;
  assign rf_MPORT_189_data = io_top_wb_bits_tc1_octet1_threadgroup4_matrix_d_data[191:128];
  assign rf_MPORT_189_addr = 8'hf7;
  assign rf_MPORT_189_mask = 1'h1;
  assign rf_MPORT_189_en = _T_162 & _GEN_15726;
  assign rf_MPORT_190_data = io_top_wb_bits_tc1_octet1_threadgroup4_matrix_d_data[127:64];
  assign rf_MPORT_190_addr = 8'hfe;
  assign rf_MPORT_190_mask = 1'h1;
  assign rf_MPORT_190_en = _T_162 & _GEN_15726;
  assign rf_MPORT_191_data = io_top_wb_bits_tc1_octet1_threadgroup4_matrix_d_data[63:0];
  assign rf_MPORT_191_addr = 8'hff;
  assign rf_MPORT_191_mask = 1'h1;
  assign rf_MPORT_191_en = _T_162 & _GEN_15726;
  assign rf_MPORT_192_data = io_uart_rf_w_data;
  assign rf_MPORT_192_addr = io_uart_rf_w_addr;
  assign rf_MPORT_192_mask = 1'h1;
  assign rf_MPORT_192_en = io_uart_rf_w_en;
  assign io_uart_ctrl_tx_en = tx_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 469:22]
  assign io_uart_rf_r_data = io_uart_rf_r_addr == 8'h0 ? 64'h0 : rf_io_uart_rf_r_data_MPORT_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 9:35]
  assign io_top_src_valid = io_top_src_valid_r; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 169:20]
  assign io_top_src_bits_tc0_ot0_tg0_matrix_a = matrix_a_0; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 176:40]
  assign io_top_src_bits_tc0_ot0_tg0_matrix_b = matrix_b_0; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 177:40]
  assign io_top_src_bits_tc0_ot0_tg0_matrix_c = matrix_c_0; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 178:40]
  assign io_top_src_bits_tc0_ot0_tg4_matrix_a = matrix_a_4; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 180:40]
  assign io_top_src_bits_tc0_ot0_tg4_matrix_b = matrix_b_4; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 181:40]
  assign io_top_src_bits_tc0_ot0_tg4_matrix_c = matrix_c_4; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 182:40]
  assign io_top_src_bits_tc0_ot1_tg0_matrix_a = matrix_a_1; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 184:40]
  assign io_top_src_bits_tc0_ot1_tg0_matrix_b = matrix_b_1; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 185:40]
  assign io_top_src_bits_tc0_ot1_tg0_matrix_c = matrix_c_1; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 186:40]
  assign io_top_src_bits_tc0_ot1_tg4_matrix_a = matrix_a_5; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 188:40]
  assign io_top_src_bits_tc0_ot1_tg4_matrix_b = matrix_b_5; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 189:40]
  assign io_top_src_bits_tc0_ot1_tg4_matrix_c = matrix_c_5; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 190:40]
  assign io_top_src_bits_tc1_ot0_tg0_matrix_a = matrix_a_2; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 192:40]
  assign io_top_src_bits_tc1_ot0_tg0_matrix_b = matrix_b_2; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 193:40]
  assign io_top_src_bits_tc1_ot0_tg0_matrix_c = matrix_c_2; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 194:40]
  assign io_top_src_bits_tc1_ot0_tg4_matrix_a = matrix_a_6; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 196:40]
  assign io_top_src_bits_tc1_ot0_tg4_matrix_b = matrix_b_6; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 197:40]
  assign io_top_src_bits_tc1_ot0_tg4_matrix_c = matrix_c_6; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 198:40]
  assign io_top_src_bits_tc1_ot1_tg0_matrix_a = matrix_a_3; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 200:40]
  assign io_top_src_bits_tc1_ot1_tg0_matrix_b = matrix_b_3; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 201:40]
  assign io_top_src_bits_tc1_ot1_tg0_matrix_c = matrix_c_3; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 202:40]
  assign io_top_src_bits_tc1_ot1_tg4_matrix_a = matrix_a_7; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 204:40]
  assign io_top_src_bits_tc1_ot1_tg4_matrix_b = matrix_b_7; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 205:40]
  assign io_top_src_bits_tc1_ot1_tg4_matrix_c = matrix_c_7; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 206:40]
  assign io_top_src_bits_ctrl_matBSel = io_top_src_bits_ctrl_mixPcMode ? step > 2'h1 : step > 2'h0; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 174:38]
  assign io_top_src_bits_ctrl_mixPcMode = io_top_src_bits_ctrl_mixPcMode_r; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 173:34]
  assign io_top_wb_ready = 1'h1; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 171:19]
  always @(posedge clock) begin
    if (rf_MPORT_en & rf_MPORT_mask) begin
      rf[rf_MPORT_addr] <= rf_MPORT_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
    end
    if (rf_MPORT_1_en & rf_MPORT_1_mask) begin
      rf[rf_MPORT_1_addr] <= rf_MPORT_1_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
    end
    if (rf_MPORT_2_en & rf_MPORT_2_mask) begin
      rf[rf_MPORT_2_addr] <= rf_MPORT_2_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
    end
    if (rf_MPORT_3_en & rf_MPORT_3_mask) begin
      rf[rf_MPORT_3_addr] <= rf_MPORT_3_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
    end
    if (rf_MPORT_4_en & rf_MPORT_4_mask) begin
      rf[rf_MPORT_4_addr] <= rf_MPORT_4_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
    end
    if (rf_MPORT_5_en & rf_MPORT_5_mask) begin
      rf[rf_MPORT_5_addr] <= rf_MPORT_5_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
    end
    if (rf_MPORT_6_en & rf_MPORT_6_mask) begin
      rf[rf_MPORT_6_addr] <= rf_MPORT_6_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
    end
    if (rf_MPORT_7_en & rf_MPORT_7_mask) begin
      rf[rf_MPORT_7_addr] <= rf_MPORT_7_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
    end
    if (rf_MPORT_8_en & rf_MPORT_8_mask) begin
      rf[rf_MPORT_8_addr] <= rf_MPORT_8_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
    end
    if (rf_MPORT_9_en & rf_MPORT_9_mask) begin
      rf[rf_MPORT_9_addr] <= rf_MPORT_9_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
    end
    if (rf_MPORT_10_en & rf_MPORT_10_mask) begin
      rf[rf_MPORT_10_addr] <= rf_MPORT_10_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
    end
    if (rf_MPORT_11_en & rf_MPORT_11_mask) begin
      rf[rf_MPORT_11_addr] <= rf_MPORT_11_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
    end
    if (rf_MPORT_12_en & rf_MPORT_12_mask) begin
      rf[rf_MPORT_12_addr] <= rf_MPORT_12_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
    end
    if (rf_MPORT_13_en & rf_MPORT_13_mask) begin
      rf[rf_MPORT_13_addr] <= rf_MPORT_13_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
    end
    if (rf_MPORT_14_en & rf_MPORT_14_mask) begin
      rf[rf_MPORT_14_addr] <= rf_MPORT_14_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
    end
    if (rf_MPORT_15_en & rf_MPORT_15_mask) begin
      rf[rf_MPORT_15_addr] <= rf_MPORT_15_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
    end
    if (rf_MPORT_16_en & rf_MPORT_16_mask) begin
      rf[rf_MPORT_16_addr] <= rf_MPORT_16_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
    end
    if (rf_MPORT_17_en & rf_MPORT_17_mask) begin
      rf[rf_MPORT_17_addr] <= rf_MPORT_17_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
    end
    if (rf_MPORT_18_en & rf_MPORT_18_mask) begin
      rf[rf_MPORT_18_addr] <= rf_MPORT_18_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
    end
    if (rf_MPORT_19_en & rf_MPORT_19_mask) begin
      rf[rf_MPORT_19_addr] <= rf_MPORT_19_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
    end
    if (rf_MPORT_20_en & rf_MPORT_20_mask) begin
      rf[rf_MPORT_20_addr] <= rf_MPORT_20_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
    end
    if (rf_MPORT_21_en & rf_MPORT_21_mask) begin
      rf[rf_MPORT_21_addr] <= rf_MPORT_21_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
    end
    if (rf_MPORT_22_en & rf_MPORT_22_mask) begin
      rf[rf_MPORT_22_addr] <= rf_MPORT_22_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
    end
    if (rf_MPORT_23_en & rf_MPORT_23_mask) begin
      rf[rf_MPORT_23_addr] <= rf_MPORT_23_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
    end
    if (rf_MPORT_24_en & rf_MPORT_24_mask) begin
      rf[rf_MPORT_24_addr] <= rf_MPORT_24_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
    end
    if (rf_MPORT_25_en & rf_MPORT_25_mask) begin
      rf[rf_MPORT_25_addr] <= rf_MPORT_25_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
    end
    if (rf_MPORT_26_en & rf_MPORT_26_mask) begin
      rf[rf_MPORT_26_addr] <= rf_MPORT_26_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
    end
    if (rf_MPORT_27_en & rf_MPORT_27_mask) begin
      rf[rf_MPORT_27_addr] <= rf_MPORT_27_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
    end
    if (rf_MPORT_28_en & rf_MPORT_28_mask) begin
      rf[rf_MPORT_28_addr] <= rf_MPORT_28_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
    end
    if (rf_MPORT_29_en & rf_MPORT_29_mask) begin
      rf[rf_MPORT_29_addr] <= rf_MPORT_29_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
    end
    if (rf_MPORT_30_en & rf_MPORT_30_mask) begin
      rf[rf_MPORT_30_addr] <= rf_MPORT_30_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
    end
    if (rf_MPORT_31_en & rf_MPORT_31_mask) begin
      rf[rf_MPORT_31_addr] <= rf_MPORT_31_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
    end
    if (rf_MPORT_32_en & rf_MPORT_32_mask) begin
      rf[rf_MPORT_32_addr] <= rf_MPORT_32_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
    end
    if (rf_MPORT_33_en & rf_MPORT_33_mask) begin
      rf[rf_MPORT_33_addr] <= rf_MPORT_33_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
    end
    if (rf_MPORT_34_en & rf_MPORT_34_mask) begin
      rf[rf_MPORT_34_addr] <= rf_MPORT_34_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
    end
    if (rf_MPORT_35_en & rf_MPORT_35_mask) begin
      rf[rf_MPORT_35_addr] <= rf_MPORT_35_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
    end
    if (rf_MPORT_36_en & rf_MPORT_36_mask) begin
      rf[rf_MPORT_36_addr] <= rf_MPORT_36_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
    end
    if (rf_MPORT_37_en & rf_MPORT_37_mask) begin
      rf[rf_MPORT_37_addr] <= rf_MPORT_37_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
    end
    if (rf_MPORT_38_en & rf_MPORT_38_mask) begin
      rf[rf_MPORT_38_addr] <= rf_MPORT_38_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
    end
    if (rf_MPORT_39_en & rf_MPORT_39_mask) begin
      rf[rf_MPORT_39_addr] <= rf_MPORT_39_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
    end
    if (rf_MPORT_40_en & rf_MPORT_40_mask) begin
      rf[rf_MPORT_40_addr] <= rf_MPORT_40_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
    end
    if (rf_MPORT_41_en & rf_MPORT_41_mask) begin
      rf[rf_MPORT_41_addr] <= rf_MPORT_41_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
    end
    if (rf_MPORT_42_en & rf_MPORT_42_mask) begin
      rf[rf_MPORT_42_addr] <= rf_MPORT_42_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
    end
    if (rf_MPORT_43_en & rf_MPORT_43_mask) begin
      rf[rf_MPORT_43_addr] <= rf_MPORT_43_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
    end
    if (rf_MPORT_44_en & rf_MPORT_44_mask) begin
      rf[rf_MPORT_44_addr] <= rf_MPORT_44_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
    end
    if (rf_MPORT_45_en & rf_MPORT_45_mask) begin
      rf[rf_MPORT_45_addr] <= rf_MPORT_45_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
    end
    if (rf_MPORT_46_en & rf_MPORT_46_mask) begin
      rf[rf_MPORT_46_addr] <= rf_MPORT_46_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
    end
    if (rf_MPORT_47_en & rf_MPORT_47_mask) begin
      rf[rf_MPORT_47_addr] <= rf_MPORT_47_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
    end
    if (rf_MPORT_48_en & rf_MPORT_48_mask) begin
      rf[rf_MPORT_48_addr] <= rf_MPORT_48_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
    end
    if (rf_MPORT_49_en & rf_MPORT_49_mask) begin
      rf[rf_MPORT_49_addr] <= rf_MPORT_49_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
    end
    if (rf_MPORT_50_en & rf_MPORT_50_mask) begin
      rf[rf_MPORT_50_addr] <= rf_MPORT_50_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
    end
    if (rf_MPORT_51_en & rf_MPORT_51_mask) begin
      rf[rf_MPORT_51_addr] <= rf_MPORT_51_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
    end
    if (rf_MPORT_52_en & rf_MPORT_52_mask) begin
      rf[rf_MPORT_52_addr] <= rf_MPORT_52_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
    end
    if (rf_MPORT_53_en & rf_MPORT_53_mask) begin
      rf[rf_MPORT_53_addr] <= rf_MPORT_53_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
    end
    if (rf_MPORT_54_en & rf_MPORT_54_mask) begin
      rf[rf_MPORT_54_addr] <= rf_MPORT_54_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
    end
    if (rf_MPORT_55_en & rf_MPORT_55_mask) begin
      rf[rf_MPORT_55_addr] <= rf_MPORT_55_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
    end
    if (rf_MPORT_56_en & rf_MPORT_56_mask) begin
      rf[rf_MPORT_56_addr] <= rf_MPORT_56_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
    end
    if (rf_MPORT_57_en & rf_MPORT_57_mask) begin
      rf[rf_MPORT_57_addr] <= rf_MPORT_57_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
    end
    if (rf_MPORT_58_en & rf_MPORT_58_mask) begin
      rf[rf_MPORT_58_addr] <= rf_MPORT_58_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
    end
    if (rf_MPORT_59_en & rf_MPORT_59_mask) begin
      rf[rf_MPORT_59_addr] <= rf_MPORT_59_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
    end
    if (rf_MPORT_60_en & rf_MPORT_60_mask) begin
      rf[rf_MPORT_60_addr] <= rf_MPORT_60_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
    end
    if (rf_MPORT_61_en & rf_MPORT_61_mask) begin
      rf[rf_MPORT_61_addr] <= rf_MPORT_61_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
    end
    if (rf_MPORT_62_en & rf_MPORT_62_mask) begin
      rf[rf_MPORT_62_addr] <= rf_MPORT_62_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
    end
    if (rf_MPORT_63_en & rf_MPORT_63_mask) begin
      rf[rf_MPORT_63_addr] <= rf_MPORT_63_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
    end
    if (rf_MPORT_64_en & rf_MPORT_64_mask) begin
      rf[rf_MPORT_64_addr] <= rf_MPORT_64_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
    end
    if (rf_MPORT_65_en & rf_MPORT_65_mask) begin
      rf[rf_MPORT_65_addr] <= rf_MPORT_65_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
    end
    if (rf_MPORT_66_en & rf_MPORT_66_mask) begin
      rf[rf_MPORT_66_addr] <= rf_MPORT_66_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
    end
    if (rf_MPORT_67_en & rf_MPORT_67_mask) begin
      rf[rf_MPORT_67_addr] <= rf_MPORT_67_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
    end
    if (rf_MPORT_68_en & rf_MPORT_68_mask) begin
      rf[rf_MPORT_68_addr] <= rf_MPORT_68_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
    end
    if (rf_MPORT_69_en & rf_MPORT_69_mask) begin
      rf[rf_MPORT_69_addr] <= rf_MPORT_69_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
    end
    if (rf_MPORT_70_en & rf_MPORT_70_mask) begin
      rf[rf_MPORT_70_addr] <= rf_MPORT_70_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
    end
    if (rf_MPORT_71_en & rf_MPORT_71_mask) begin
      rf[rf_MPORT_71_addr] <= rf_MPORT_71_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
    end
    if (rf_MPORT_72_en & rf_MPORT_72_mask) begin
      rf[rf_MPORT_72_addr] <= rf_MPORT_72_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
    end
    if (rf_MPORT_73_en & rf_MPORT_73_mask) begin
      rf[rf_MPORT_73_addr] <= rf_MPORT_73_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
    end
    if (rf_MPORT_74_en & rf_MPORT_74_mask) begin
      rf[rf_MPORT_74_addr] <= rf_MPORT_74_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
    end
    if (rf_MPORT_75_en & rf_MPORT_75_mask) begin
      rf[rf_MPORT_75_addr] <= rf_MPORT_75_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
    end
    if (rf_MPORT_76_en & rf_MPORT_76_mask) begin
      rf[rf_MPORT_76_addr] <= rf_MPORT_76_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
    end
    if (rf_MPORT_77_en & rf_MPORT_77_mask) begin
      rf[rf_MPORT_77_addr] <= rf_MPORT_77_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
    end
    if (rf_MPORT_78_en & rf_MPORT_78_mask) begin
      rf[rf_MPORT_78_addr] <= rf_MPORT_78_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
    end
    if (rf_MPORT_79_en & rf_MPORT_79_mask) begin
      rf[rf_MPORT_79_addr] <= rf_MPORT_79_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
    end
    if (rf_MPORT_80_en & rf_MPORT_80_mask) begin
      rf[rf_MPORT_80_addr] <= rf_MPORT_80_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
    end
    if (rf_MPORT_81_en & rf_MPORT_81_mask) begin
      rf[rf_MPORT_81_addr] <= rf_MPORT_81_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
    end
    if (rf_MPORT_82_en & rf_MPORT_82_mask) begin
      rf[rf_MPORT_82_addr] <= rf_MPORT_82_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
    end
    if (rf_MPORT_83_en & rf_MPORT_83_mask) begin
      rf[rf_MPORT_83_addr] <= rf_MPORT_83_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
    end
    if (rf_MPORT_84_en & rf_MPORT_84_mask) begin
      rf[rf_MPORT_84_addr] <= rf_MPORT_84_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
    end
    if (rf_MPORT_85_en & rf_MPORT_85_mask) begin
      rf[rf_MPORT_85_addr] <= rf_MPORT_85_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
    end
    if (rf_MPORT_86_en & rf_MPORT_86_mask) begin
      rf[rf_MPORT_86_addr] <= rf_MPORT_86_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
    end
    if (rf_MPORT_87_en & rf_MPORT_87_mask) begin
      rf[rf_MPORT_87_addr] <= rf_MPORT_87_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
    end
    if (rf_MPORT_88_en & rf_MPORT_88_mask) begin
      rf[rf_MPORT_88_addr] <= rf_MPORT_88_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
    end
    if (rf_MPORT_89_en & rf_MPORT_89_mask) begin
      rf[rf_MPORT_89_addr] <= rf_MPORT_89_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
    end
    if (rf_MPORT_90_en & rf_MPORT_90_mask) begin
      rf[rf_MPORT_90_addr] <= rf_MPORT_90_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
    end
    if (rf_MPORT_91_en & rf_MPORT_91_mask) begin
      rf[rf_MPORT_91_addr] <= rf_MPORT_91_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
    end
    if (rf_MPORT_92_en & rf_MPORT_92_mask) begin
      rf[rf_MPORT_92_addr] <= rf_MPORT_92_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
    end
    if (rf_MPORT_93_en & rf_MPORT_93_mask) begin
      rf[rf_MPORT_93_addr] <= rf_MPORT_93_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
    end
    if (rf_MPORT_94_en & rf_MPORT_94_mask) begin
      rf[rf_MPORT_94_addr] <= rf_MPORT_94_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
    end
    if (rf_MPORT_95_en & rf_MPORT_95_mask) begin
      rf[rf_MPORT_95_addr] <= rf_MPORT_95_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
    end
    if (rf_MPORT_96_en & rf_MPORT_96_mask) begin
      rf[rf_MPORT_96_addr] <= rf_MPORT_96_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
    end
    if (rf_MPORT_97_en & rf_MPORT_97_mask) begin
      rf[rf_MPORT_97_addr] <= rf_MPORT_97_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
    end
    if (rf_MPORT_98_en & rf_MPORT_98_mask) begin
      rf[rf_MPORT_98_addr] <= rf_MPORT_98_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
    end
    if (rf_MPORT_99_en & rf_MPORT_99_mask) begin
      rf[rf_MPORT_99_addr] <= rf_MPORT_99_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
    end
    if (rf_MPORT_100_en & rf_MPORT_100_mask) begin
      rf[rf_MPORT_100_addr] <= rf_MPORT_100_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
    end
    if (rf_MPORT_101_en & rf_MPORT_101_mask) begin
      rf[rf_MPORT_101_addr] <= rf_MPORT_101_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
    end
    if (rf_MPORT_102_en & rf_MPORT_102_mask) begin
      rf[rf_MPORT_102_addr] <= rf_MPORT_102_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
    end
    if (rf_MPORT_103_en & rf_MPORT_103_mask) begin
      rf[rf_MPORT_103_addr] <= rf_MPORT_103_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
    end
    if (rf_MPORT_104_en & rf_MPORT_104_mask) begin
      rf[rf_MPORT_104_addr] <= rf_MPORT_104_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
    end
    if (rf_MPORT_105_en & rf_MPORT_105_mask) begin
      rf[rf_MPORT_105_addr] <= rf_MPORT_105_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
    end
    if (rf_MPORT_106_en & rf_MPORT_106_mask) begin
      rf[rf_MPORT_106_addr] <= rf_MPORT_106_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
    end
    if (rf_MPORT_107_en & rf_MPORT_107_mask) begin
      rf[rf_MPORT_107_addr] <= rf_MPORT_107_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
    end
    if (rf_MPORT_108_en & rf_MPORT_108_mask) begin
      rf[rf_MPORT_108_addr] <= rf_MPORT_108_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
    end
    if (rf_MPORT_109_en & rf_MPORT_109_mask) begin
      rf[rf_MPORT_109_addr] <= rf_MPORT_109_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
    end
    if (rf_MPORT_110_en & rf_MPORT_110_mask) begin
      rf[rf_MPORT_110_addr] <= rf_MPORT_110_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
    end
    if (rf_MPORT_111_en & rf_MPORT_111_mask) begin
      rf[rf_MPORT_111_addr] <= rf_MPORT_111_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
    end
    if (rf_MPORT_112_en & rf_MPORT_112_mask) begin
      rf[rf_MPORT_112_addr] <= rf_MPORT_112_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
    end
    if (rf_MPORT_113_en & rf_MPORT_113_mask) begin
      rf[rf_MPORT_113_addr] <= rf_MPORT_113_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
    end
    if (rf_MPORT_114_en & rf_MPORT_114_mask) begin
      rf[rf_MPORT_114_addr] <= rf_MPORT_114_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
    end
    if (rf_MPORT_115_en & rf_MPORT_115_mask) begin
      rf[rf_MPORT_115_addr] <= rf_MPORT_115_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
    end
    if (rf_MPORT_116_en & rf_MPORT_116_mask) begin
      rf[rf_MPORT_116_addr] <= rf_MPORT_116_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
    end
    if (rf_MPORT_117_en & rf_MPORT_117_mask) begin
      rf[rf_MPORT_117_addr] <= rf_MPORT_117_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
    end
    if (rf_MPORT_118_en & rf_MPORT_118_mask) begin
      rf[rf_MPORT_118_addr] <= rf_MPORT_118_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
    end
    if (rf_MPORT_119_en & rf_MPORT_119_mask) begin
      rf[rf_MPORT_119_addr] <= rf_MPORT_119_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
    end
    if (rf_MPORT_120_en & rf_MPORT_120_mask) begin
      rf[rf_MPORT_120_addr] <= rf_MPORT_120_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
    end
    if (rf_MPORT_121_en & rf_MPORT_121_mask) begin
      rf[rf_MPORT_121_addr] <= rf_MPORT_121_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
    end
    if (rf_MPORT_122_en & rf_MPORT_122_mask) begin
      rf[rf_MPORT_122_addr] <= rf_MPORT_122_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
    end
    if (rf_MPORT_123_en & rf_MPORT_123_mask) begin
      rf[rf_MPORT_123_addr] <= rf_MPORT_123_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
    end
    if (rf_MPORT_124_en & rf_MPORT_124_mask) begin
      rf[rf_MPORT_124_addr] <= rf_MPORT_124_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
    end
    if (rf_MPORT_125_en & rf_MPORT_125_mask) begin
      rf[rf_MPORT_125_addr] <= rf_MPORT_125_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
    end
    if (rf_MPORT_126_en & rf_MPORT_126_mask) begin
      rf[rf_MPORT_126_addr] <= rf_MPORT_126_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
    end
    if (rf_MPORT_127_en & rf_MPORT_127_mask) begin
      rf[rf_MPORT_127_addr] <= rf_MPORT_127_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
    end
    if (rf_MPORT_128_en & rf_MPORT_128_mask) begin
      rf[rf_MPORT_128_addr] <= rf_MPORT_128_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
    end
    if (rf_MPORT_129_en & rf_MPORT_129_mask) begin
      rf[rf_MPORT_129_addr] <= rf_MPORT_129_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
    end
    if (rf_MPORT_130_en & rf_MPORT_130_mask) begin
      rf[rf_MPORT_130_addr] <= rf_MPORT_130_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
    end
    if (rf_MPORT_131_en & rf_MPORT_131_mask) begin
      rf[rf_MPORT_131_addr] <= rf_MPORT_131_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
    end
    if (rf_MPORT_132_en & rf_MPORT_132_mask) begin
      rf[rf_MPORT_132_addr] <= rf_MPORT_132_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
    end
    if (rf_MPORT_133_en & rf_MPORT_133_mask) begin
      rf[rf_MPORT_133_addr] <= rf_MPORT_133_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
    end
    if (rf_MPORT_134_en & rf_MPORT_134_mask) begin
      rf[rf_MPORT_134_addr] <= rf_MPORT_134_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
    end
    if (rf_MPORT_135_en & rf_MPORT_135_mask) begin
      rf[rf_MPORT_135_addr] <= rf_MPORT_135_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
    end
    if (rf_MPORT_136_en & rf_MPORT_136_mask) begin
      rf[rf_MPORT_136_addr] <= rf_MPORT_136_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
    end
    if (rf_MPORT_137_en & rf_MPORT_137_mask) begin
      rf[rf_MPORT_137_addr] <= rf_MPORT_137_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
    end
    if (rf_MPORT_138_en & rf_MPORT_138_mask) begin
      rf[rf_MPORT_138_addr] <= rf_MPORT_138_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
    end
    if (rf_MPORT_139_en & rf_MPORT_139_mask) begin
      rf[rf_MPORT_139_addr] <= rf_MPORT_139_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
    end
    if (rf_MPORT_140_en & rf_MPORT_140_mask) begin
      rf[rf_MPORT_140_addr] <= rf_MPORT_140_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
    end
    if (rf_MPORT_141_en & rf_MPORT_141_mask) begin
      rf[rf_MPORT_141_addr] <= rf_MPORT_141_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
    end
    if (rf_MPORT_142_en & rf_MPORT_142_mask) begin
      rf[rf_MPORT_142_addr] <= rf_MPORT_142_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
    end
    if (rf_MPORT_143_en & rf_MPORT_143_mask) begin
      rf[rf_MPORT_143_addr] <= rf_MPORT_143_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
    end
    if (rf_MPORT_144_en & rf_MPORT_144_mask) begin
      rf[rf_MPORT_144_addr] <= rf_MPORT_144_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
    end
    if (rf_MPORT_145_en & rf_MPORT_145_mask) begin
      rf[rf_MPORT_145_addr] <= rf_MPORT_145_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
    end
    if (rf_MPORT_146_en & rf_MPORT_146_mask) begin
      rf[rf_MPORT_146_addr] <= rf_MPORT_146_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
    end
    if (rf_MPORT_147_en & rf_MPORT_147_mask) begin
      rf[rf_MPORT_147_addr] <= rf_MPORT_147_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
    end
    if (rf_MPORT_148_en & rf_MPORT_148_mask) begin
      rf[rf_MPORT_148_addr] <= rf_MPORT_148_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
    end
    if (rf_MPORT_149_en & rf_MPORT_149_mask) begin
      rf[rf_MPORT_149_addr] <= rf_MPORT_149_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
    end
    if (rf_MPORT_150_en & rf_MPORT_150_mask) begin
      rf[rf_MPORT_150_addr] <= rf_MPORT_150_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
    end
    if (rf_MPORT_151_en & rf_MPORT_151_mask) begin
      rf[rf_MPORT_151_addr] <= rf_MPORT_151_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
    end
    if (rf_MPORT_152_en & rf_MPORT_152_mask) begin
      rf[rf_MPORT_152_addr] <= rf_MPORT_152_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
    end
    if (rf_MPORT_153_en & rf_MPORT_153_mask) begin
      rf[rf_MPORT_153_addr] <= rf_MPORT_153_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
    end
    if (rf_MPORT_154_en & rf_MPORT_154_mask) begin
      rf[rf_MPORT_154_addr] <= rf_MPORT_154_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
    end
    if (rf_MPORT_155_en & rf_MPORT_155_mask) begin
      rf[rf_MPORT_155_addr] <= rf_MPORT_155_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
    end
    if (rf_MPORT_156_en & rf_MPORT_156_mask) begin
      rf[rf_MPORT_156_addr] <= rf_MPORT_156_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
    end
    if (rf_MPORT_157_en & rf_MPORT_157_mask) begin
      rf[rf_MPORT_157_addr] <= rf_MPORT_157_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
    end
    if (rf_MPORT_158_en & rf_MPORT_158_mask) begin
      rf[rf_MPORT_158_addr] <= rf_MPORT_158_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
    end
    if (rf_MPORT_159_en & rf_MPORT_159_mask) begin
      rf[rf_MPORT_159_addr] <= rf_MPORT_159_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
    end
    if (rf_MPORT_160_en & rf_MPORT_160_mask) begin
      rf[rf_MPORT_160_addr] <= rf_MPORT_160_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
    end
    if (rf_MPORT_161_en & rf_MPORT_161_mask) begin
      rf[rf_MPORT_161_addr] <= rf_MPORT_161_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
    end
    if (rf_MPORT_162_en & rf_MPORT_162_mask) begin
      rf[rf_MPORT_162_addr] <= rf_MPORT_162_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
    end
    if (rf_MPORT_163_en & rf_MPORT_163_mask) begin
      rf[rf_MPORT_163_addr] <= rf_MPORT_163_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
    end
    if (rf_MPORT_164_en & rf_MPORT_164_mask) begin
      rf[rf_MPORT_164_addr] <= rf_MPORT_164_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
    end
    if (rf_MPORT_165_en & rf_MPORT_165_mask) begin
      rf[rf_MPORT_165_addr] <= rf_MPORT_165_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
    end
    if (rf_MPORT_166_en & rf_MPORT_166_mask) begin
      rf[rf_MPORT_166_addr] <= rf_MPORT_166_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
    end
    if (rf_MPORT_167_en & rf_MPORT_167_mask) begin
      rf[rf_MPORT_167_addr] <= rf_MPORT_167_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
    end
    if (rf_MPORT_168_en & rf_MPORT_168_mask) begin
      rf[rf_MPORT_168_addr] <= rf_MPORT_168_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
    end
    if (rf_MPORT_169_en & rf_MPORT_169_mask) begin
      rf[rf_MPORT_169_addr] <= rf_MPORT_169_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
    end
    if (rf_MPORT_170_en & rf_MPORT_170_mask) begin
      rf[rf_MPORT_170_addr] <= rf_MPORT_170_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
    end
    if (rf_MPORT_171_en & rf_MPORT_171_mask) begin
      rf[rf_MPORT_171_addr] <= rf_MPORT_171_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
    end
    if (rf_MPORT_172_en & rf_MPORT_172_mask) begin
      rf[rf_MPORT_172_addr] <= rf_MPORT_172_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
    end
    if (rf_MPORT_173_en & rf_MPORT_173_mask) begin
      rf[rf_MPORT_173_addr] <= rf_MPORT_173_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
    end
    if (rf_MPORT_174_en & rf_MPORT_174_mask) begin
      rf[rf_MPORT_174_addr] <= rf_MPORT_174_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
    end
    if (rf_MPORT_175_en & rf_MPORT_175_mask) begin
      rf[rf_MPORT_175_addr] <= rf_MPORT_175_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
    end
    if (rf_MPORT_176_en & rf_MPORT_176_mask) begin
      rf[rf_MPORT_176_addr] <= rf_MPORT_176_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
    end
    if (rf_MPORT_177_en & rf_MPORT_177_mask) begin
      rf[rf_MPORT_177_addr] <= rf_MPORT_177_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
    end
    if (rf_MPORT_178_en & rf_MPORT_178_mask) begin
      rf[rf_MPORT_178_addr] <= rf_MPORT_178_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
    end
    if (rf_MPORT_179_en & rf_MPORT_179_mask) begin
      rf[rf_MPORT_179_addr] <= rf_MPORT_179_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
    end
    if (rf_MPORT_180_en & rf_MPORT_180_mask) begin
      rf[rf_MPORT_180_addr] <= rf_MPORT_180_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
    end
    if (rf_MPORT_181_en & rf_MPORT_181_mask) begin
      rf[rf_MPORT_181_addr] <= rf_MPORT_181_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
    end
    if (rf_MPORT_182_en & rf_MPORT_182_mask) begin
      rf[rf_MPORT_182_addr] <= rf_MPORT_182_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
    end
    if (rf_MPORT_183_en & rf_MPORT_183_mask) begin
      rf[rf_MPORT_183_addr] <= rf_MPORT_183_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
    end
    if (rf_MPORT_184_en & rf_MPORT_184_mask) begin
      rf[rf_MPORT_184_addr] <= rf_MPORT_184_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
    end
    if (rf_MPORT_185_en & rf_MPORT_185_mask) begin
      rf[rf_MPORT_185_addr] <= rf_MPORT_185_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
    end
    if (rf_MPORT_186_en & rf_MPORT_186_mask) begin
      rf[rf_MPORT_186_addr] <= rf_MPORT_186_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
    end
    if (rf_MPORT_187_en & rf_MPORT_187_mask) begin
      rf[rf_MPORT_187_addr] <= rf_MPORT_187_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
    end
    if (rf_MPORT_188_en & rf_MPORT_188_mask) begin
      rf[rf_MPORT_188_addr] <= rf_MPORT_188_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
    end
    if (rf_MPORT_189_en & rf_MPORT_189_mask) begin
      rf[rf_MPORT_189_addr] <= rf_MPORT_189_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
    end
    if (rf_MPORT_190_en & rf_MPORT_190_mask) begin
      rf[rf_MPORT_190_addr] <= rf_MPORT_190_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
    end
    if (rf_MPORT_191_en & rf_MPORT_191_mask) begin
      rf[rf_MPORT_191_addr] <= rf_MPORT_191_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
    end
    if (rf_MPORT_192_en & rf_MPORT_192_mask) begin
      rf[rf_MPORT_192_addr] <= rf_MPORT_192_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 8:15]
    end
    if (reset) begin // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 146:20]
      set <= 2'h0; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 146:20]
    end else if (handshaked) begin // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 208:20]
      if (step == MAX_STEP) begin // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 382:29]
        set <= _set_T_1; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 387:11]
      end
    end
    if (reset) begin // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 147:21]
      step <= 2'h0; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 147:21]
    end else if (handshaked) begin // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 208:20]
      if (step == MAX_STEP) begin // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 382:29]
        step <= 2'h0; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 383:12]
      end else begin
        step <= _step_T_1; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 389:12]
      end
    end
    if (reset) begin // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 148:24]
      out_set <= 2'h0; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 148:24]
    end else if (_T_162) begin // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 393:24]
      if (out_step == MAX_STEP) begin // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 459:33]
        out_set <= _out_set_T_1; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 464:15]
      end
    end
    if (reset) begin // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 149:25]
      out_step <= 2'h0; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 149:25]
    end else if (_T_162) begin // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 393:24]
      if (out_step == MAX_STEP) begin // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 459:33]
        out_step <= 2'h0; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 460:16]
      end else begin
        out_step <= _out_step_T_1; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 466:16]
      end
    end
    if (reset) begin // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 150:24]
      exec_en <= 1'h0; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 150:24]
    end else if (handshaked) begin // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 208:20]
      if (step == MAX_STEP) begin // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 382:29]
        if (set == 2'h3) begin // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 384:34]
          exec_en <= 1'h0; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 385:17]
        end else begin
          exec_en <= _GEN_0;
        end
      end else begin
        exec_en <= _GEN_0;
      end
    end else begin
      exec_en <= _GEN_0;
    end
    if (reset) begin // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 154:22]
      tx_en <= 1'h0; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 154:22]
    end else if (_T_162) begin // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 393:24]
      if (out_step == MAX_STEP) begin // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 459:33]
        tx_en <= _GEN_15791;
      end else begin
        tx_en <= _GEN_1;
      end
    end else begin
      tx_en <= _GEN_1;
    end
    if (handshaked) begin // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 208:20]
      if (2'h0 == set) begin // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 210:18]
        if (2'h0 == step) begin // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 212:23]
          if (io_mixPc) begin // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 214:29]
            matrix_a_0 <= _matrix_a_0_T; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 216:29]
          end else begin
            matrix_a_0 <= a_1; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 221:29]
          end
        end else if (2'h1 == step) begin // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 212:23]
          matrix_a_0 <= _GEN_36;
        end else begin
          matrix_a_0 <= _GEN_66;
        end
      end else if (2'h1 == set) begin // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 210:18]
        if (_T_1) begin // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 254:24]
          matrix_a_0 <= _GEN_223;
        end else begin
          matrix_a_0 <= _GEN_289;
        end
      end else if (2'h2 == set) begin // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 210:18]
        matrix_a_0 <= _GEN_538;
      end else begin
        matrix_a_0 <= _GEN_813;
      end
    end
    if (handshaked) begin // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 208:20]
      if (2'h0 == set) begin // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 210:18]
        if (2'h0 == step) begin // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 212:23]
          if (io_mixPc) begin // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 214:29]
            matrix_a_1 <= _matrix_a_1_T; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 216:29]
          end else begin
            matrix_a_1 <= a_25; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 221:29]
          end
        end else if (2'h1 == step) begin // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 212:23]
          matrix_a_1 <= _GEN_1600;
        end else begin
          matrix_a_1 <= _GEN_1630;
        end
      end else if (2'h1 == set) begin // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 210:18]
        if (_T_1) begin // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 254:24]
          matrix_a_1 <= _GEN_1787;
        end else begin
          matrix_a_1 <= _GEN_1845;
        end
      end else if (2'h2 == set) begin // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 210:18]
        matrix_a_1 <= _GEN_2086;
      end else begin
        matrix_a_1 <= _GEN_2353;
      end
    end
    if (handshaked) begin // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 208:20]
      if (2'h0 == set) begin // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 210:18]
        if (2'h0 == step) begin // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 212:23]
          if (io_mixPc) begin // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 214:29]
            matrix_a_2 <= _matrix_a_2_T; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 216:29]
          end else begin
            matrix_a_2 <= a_49; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 221:29]
          end
        end else if (2'h1 == step) begin // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 212:23]
          matrix_a_2 <= _GEN_3140;
        end else begin
          matrix_a_2 <= _GEN_3170;
        end
      end else if (2'h1 == set) begin // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 210:18]
        if (_T_1) begin // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 254:24]
          matrix_a_2 <= _GEN_3325;
        end else begin
          matrix_a_2 <= _GEN_3385;
        end
      end else if (2'h2 == set) begin // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 210:18]
        matrix_a_2 <= _GEN_3626;
      end else begin
        matrix_a_2 <= _GEN_3893;
      end
    end
    if (handshaked) begin // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 208:20]
      if (2'h0 == set) begin // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 210:18]
        if (2'h0 == step) begin // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 212:23]
          if (io_mixPc) begin // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 214:29]
            matrix_a_3 <= _matrix_a_3_T; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 216:29]
          end else begin
            matrix_a_3 <= a_73; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 221:29]
          end
        end else if (2'h1 == step) begin // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 212:23]
          matrix_a_3 <= _GEN_4672;
        end else begin
          matrix_a_3 <= _GEN_4702;
        end
      end else if (2'h1 == set) begin // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 210:18]
        if (_T_1) begin // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 254:24]
          matrix_a_3 <= _GEN_4857;
        end else begin
          matrix_a_3 <= _GEN_4909;
        end
      end else if (2'h2 == set) begin // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 210:18]
        matrix_a_3 <= _GEN_5142;
      end else begin
        matrix_a_3 <= _GEN_5401;
      end
    end
    if (handshaked) begin // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 208:20]
      if (2'h0 == set) begin // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 210:18]
        if (2'h0 == step) begin // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 212:23]
          if (io_mixPc) begin // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 214:29]
            matrix_a_4 <= _matrix_a_4_T; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 216:29]
          end else begin
            matrix_a_4 <= a_97; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 221:29]
          end
        end else if (2'h1 == step) begin // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 212:23]
          matrix_a_4 <= _GEN_6196;
        end else begin
          matrix_a_4 <= _GEN_6226;
        end
      end else if (2'h1 == set) begin // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 210:18]
        if (_T_1) begin // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 254:24]
          matrix_a_4 <= _GEN_6383;
        end else begin
          matrix_a_4 <= _GEN_6449;
        end
      end else if (2'h2 == set) begin // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 210:18]
        matrix_a_4 <= _GEN_6698;
      end else begin
        matrix_a_4 <= _GEN_6973;
      end
    end
    if (handshaked) begin // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 208:20]
      if (2'h0 == set) begin // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 210:18]
        if (2'h0 == step) begin // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 212:23]
          if (io_mixPc) begin // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 214:29]
            matrix_a_5 <= _matrix_a_5_T; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 216:29]
          end else begin
            matrix_a_5 <= a_121; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 221:29]
          end
        end else if (2'h1 == step) begin // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 212:23]
          matrix_a_5 <= _GEN_7760;
        end else begin
          matrix_a_5 <= _GEN_7790;
        end
      end else if (2'h1 == set) begin // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 210:18]
        if (_T_1) begin // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 254:24]
          matrix_a_5 <= _GEN_7947;
        end else begin
          matrix_a_5 <= _GEN_8005;
        end
      end else if (2'h2 == set) begin // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 210:18]
        matrix_a_5 <= _GEN_8246;
      end else begin
        matrix_a_5 <= _GEN_8513;
      end
    end
    if (handshaked) begin // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 208:20]
      if (2'h0 == set) begin // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 210:18]
        if (2'h0 == step) begin // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 212:23]
          if (io_mixPc) begin // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 214:29]
            matrix_a_6 <= _matrix_a_6_T; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 216:29]
          end else begin
            matrix_a_6 <= a_145; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 221:29]
          end
        end else if (2'h1 == step) begin // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 212:23]
          matrix_a_6 <= _GEN_9300;
        end else begin
          matrix_a_6 <= _GEN_9330;
        end
      end else if (2'h1 == set) begin // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 210:18]
        if (_T_1) begin // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 254:24]
          matrix_a_6 <= _GEN_9485;
        end else begin
          matrix_a_6 <= _GEN_9545;
        end
      end else if (2'h2 == set) begin // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 210:18]
        matrix_a_6 <= _GEN_9786;
      end else begin
        matrix_a_6 <= _GEN_10053;
      end
    end
    if (handshaked) begin // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 208:20]
      if (2'h0 == set) begin // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 210:18]
        if (2'h0 == step) begin // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 212:23]
          if (io_mixPc) begin // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 214:29]
            matrix_a_7 <= _matrix_a_7_T; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 216:29]
          end else begin
            matrix_a_7 <= a_169; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 221:29]
          end
        end else if (2'h1 == step) begin // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 212:23]
          matrix_a_7 <= _GEN_10832;
        end else begin
          matrix_a_7 <= _GEN_10862;
        end
      end else if (2'h1 == set) begin // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 210:18]
        if (_T_1) begin // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 254:24]
          matrix_a_7 <= _GEN_11017;
        end else begin
          matrix_a_7 <= _GEN_11069;
        end
      end else if (2'h2 == set) begin // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 210:18]
        matrix_a_7 <= _GEN_11302;
      end else begin
        matrix_a_7 <= _GEN_11561;
      end
    end
    if (handshaked) begin // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 208:20]
      if (2'h0 == set) begin // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 210:18]
        if (2'h0 == step) begin // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 212:23]
          if (io_mixPc) begin // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 214:29]
            matrix_b_0 <= _matrix_b_0_T; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 217:29]
          end else begin
            matrix_b_0 <= _matrix_b_0_T_1; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 222:29]
          end
        end else if (2'h1 == step) begin // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 212:23]
          matrix_b_0 <= _GEN_37;
        end else begin
          matrix_b_0 <= _GEN_71;
        end
      end else if (2'h1 == set) begin // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 210:18]
        if (_T_1) begin // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 254:24]
          matrix_b_0 <= _GEN_228;
        end else begin
          matrix_b_0 <= _GEN_294;
        end
      end else if (2'h2 == set) begin // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 210:18]
        matrix_b_0 <= _GEN_543;
      end else begin
        matrix_b_0 <= _GEN_818;
      end
    end
    if (handshaked) begin // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 208:20]
      if (2'h0 == set) begin // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 210:18]
        if (2'h0 == step) begin // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 212:23]
          if (io_mixPc) begin // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 214:29]
            matrix_b_1 <= _matrix_b_1_T; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 217:29]
          end else begin
            matrix_b_1 <= _matrix_b_1_T_1; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 222:29]
          end
        end else if (2'h1 == step) begin // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 212:23]
          matrix_b_1 <= _GEN_1601;
        end else begin
          matrix_b_1 <= _GEN_1635;
        end
      end else if (2'h1 == set) begin // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 210:18]
        if (_T_1) begin // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 254:24]
          matrix_b_1 <= _GEN_1788;
        end else begin
          matrix_b_1 <= _GEN_1850;
        end
      end else if (2'h2 == set) begin // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 210:18]
        matrix_b_1 <= _GEN_2091;
      end else begin
        matrix_b_1 <= _GEN_2358;
      end
    end
    if (handshaked) begin // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 208:20]
      if (2'h0 == set) begin // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 210:18]
        if (2'h0 == step) begin // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 212:23]
          if (io_mixPc) begin // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 214:29]
            matrix_b_2 <= _matrix_b_2_T; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 217:29]
          end else begin
            matrix_b_2 <= _matrix_b_2_T_1; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 222:29]
          end
        end else if (2'h1 == step) begin // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 212:23]
          matrix_b_2 <= _GEN_3141;
        end else begin
          matrix_b_2 <= _GEN_3175;
        end
      end else if (2'h1 == set) begin // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 210:18]
        if (_T_1) begin // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 254:24]
          matrix_b_2 <= _GEN_3330;
        end else begin
          matrix_b_2 <= _GEN_3390;
        end
      end else if (2'h2 == set) begin // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 210:18]
        matrix_b_2 <= _GEN_3631;
      end else begin
        matrix_b_2 <= _GEN_3898;
      end
    end
    if (handshaked) begin // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 208:20]
      if (2'h0 == set) begin // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 210:18]
        if (2'h0 == step) begin // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 212:23]
          if (io_mixPc) begin // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 214:29]
            matrix_b_3 <= _matrix_b_3_T; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 217:29]
          end else begin
            matrix_b_3 <= _matrix_b_3_T_1; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 222:29]
          end
        end else if (2'h1 == step) begin // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 212:23]
          matrix_b_3 <= _GEN_4673;
        end else begin
          matrix_b_3 <= _GEN_4707;
        end
      end else if (2'h1 == set) begin // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 210:18]
        if (_T_1) begin // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 254:24]
          matrix_b_3 <= _GEN_4858;
        end else begin
          matrix_b_3 <= _GEN_4914;
        end
      end else if (2'h2 == set) begin // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 210:18]
        matrix_b_3 <= _GEN_5147;
      end else begin
        matrix_b_3 <= _GEN_5406;
      end
    end
    if (handshaked) begin // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 208:20]
      if (2'h0 == set) begin // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 210:18]
        if (2'h0 == step) begin // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 212:23]
          if (io_mixPc) begin // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 214:29]
            matrix_b_4 <= _matrix_b_4_T; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 217:29]
          end else begin
            matrix_b_4 <= _matrix_b_4_T_1; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 222:29]
          end
        end else if (2'h1 == step) begin // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 212:23]
          matrix_b_4 <= _GEN_6197;
        end else begin
          matrix_b_4 <= _GEN_6231;
        end
      end else if (2'h1 == set) begin // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 210:18]
        if (_T_1) begin // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 254:24]
          matrix_b_4 <= _GEN_6388;
        end else begin
          matrix_b_4 <= _GEN_6454;
        end
      end else if (2'h2 == set) begin // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 210:18]
        matrix_b_4 <= _GEN_6703;
      end else begin
        matrix_b_4 <= _GEN_6978;
      end
    end
    if (handshaked) begin // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 208:20]
      if (2'h0 == set) begin // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 210:18]
        if (2'h0 == step) begin // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 212:23]
          if (io_mixPc) begin // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 214:29]
            matrix_b_5 <= _matrix_b_5_T; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 217:29]
          end else begin
            matrix_b_5 <= _matrix_b_5_T_1; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 222:29]
          end
        end else if (2'h1 == step) begin // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 212:23]
          matrix_b_5 <= _GEN_7761;
        end else begin
          matrix_b_5 <= _GEN_7795;
        end
      end else if (2'h1 == set) begin // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 210:18]
        if (_T_1) begin // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 254:24]
          matrix_b_5 <= _GEN_7948;
        end else begin
          matrix_b_5 <= _GEN_8010;
        end
      end else if (2'h2 == set) begin // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 210:18]
        matrix_b_5 <= _GEN_8251;
      end else begin
        matrix_b_5 <= _GEN_8518;
      end
    end
    if (handshaked) begin // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 208:20]
      if (2'h0 == set) begin // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 210:18]
        if (2'h0 == step) begin // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 212:23]
          if (io_mixPc) begin // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 214:29]
            matrix_b_6 <= _matrix_b_6_T; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 217:29]
          end else begin
            matrix_b_6 <= _matrix_b_6_T_1; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 222:29]
          end
        end else if (2'h1 == step) begin // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 212:23]
          matrix_b_6 <= _GEN_9301;
        end else begin
          matrix_b_6 <= _GEN_9335;
        end
      end else if (2'h1 == set) begin // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 210:18]
        if (_T_1) begin // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 254:24]
          matrix_b_6 <= _GEN_9490;
        end else begin
          matrix_b_6 <= _GEN_9550;
        end
      end else if (2'h2 == set) begin // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 210:18]
        matrix_b_6 <= _GEN_9791;
      end else begin
        matrix_b_6 <= _GEN_10058;
      end
    end
    if (handshaked) begin // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 208:20]
      if (2'h0 == set) begin // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 210:18]
        if (2'h0 == step) begin // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 212:23]
          if (io_mixPc) begin // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 214:29]
            matrix_b_7 <= _matrix_b_7_T; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 217:29]
          end else begin
            matrix_b_7 <= _matrix_b_7_T_1; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 222:29]
          end
        end else if (2'h1 == step) begin // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 212:23]
          matrix_b_7 <= _GEN_10833;
        end else begin
          matrix_b_7 <= _GEN_10867;
        end
      end else if (2'h1 == set) begin // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 210:18]
        if (_T_1) begin // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 254:24]
          matrix_b_7 <= _GEN_11018;
        end else begin
          matrix_b_7 <= _GEN_11074;
        end
      end else if (2'h2 == set) begin // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 210:18]
        matrix_b_7 <= _GEN_11307;
      end else begin
        matrix_b_7 <= _GEN_11566;
      end
    end
    if (handshaked) begin // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 208:20]
      if (2'h0 == set) begin // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 210:18]
        if (2'h0 == step) begin // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 212:23]
          if (io_mixPc) begin // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 214:29]
            matrix_c_0 <= _matrix_c_0_T; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 218:29]
          end else begin
            matrix_c_0 <= _matrix_c_0_T_1; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 223:29]
          end
        end else if (2'h1 == step) begin // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 212:23]
          matrix_c_0 <= _GEN_42;
        end else begin
          matrix_c_0 <= _GEN_76;
        end
      end else if (2'h1 == set) begin // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 210:18]
        if (_T_1) begin // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 254:24]
          matrix_c_0 <= _GEN_229;
        end else begin
          matrix_c_0 <= _GEN_299;
        end
      end else if (2'h2 == set) begin // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 210:18]
        matrix_c_0 <= _GEN_548;
      end else begin
        matrix_c_0 <= _GEN_823;
      end
    end
    if (handshaked) begin // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 208:20]
      if (2'h0 == set) begin // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 210:18]
        if (2'h0 == step) begin // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 212:23]
          if (io_mixPc) begin // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 214:29]
            matrix_c_1 <= _matrix_c_1_T; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 218:29]
          end else begin
            matrix_c_1 <= _matrix_c_1_T_1; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 223:29]
          end
        end else if (2'h1 == step) begin // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 212:23]
          matrix_c_1 <= _GEN_1606;
        end else begin
          matrix_c_1 <= _GEN_1640;
        end
      end else if (2'h1 == set) begin // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 210:18]
        if (_T_1) begin // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 254:24]
          matrix_c_1 <= _GEN_1789;
        end else begin
          matrix_c_1 <= _GEN_1855;
        end
      end else if (2'h2 == set) begin // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 210:18]
        matrix_c_1 <= _GEN_2096;
      end else begin
        matrix_c_1 <= _GEN_2363;
      end
    end
    if (handshaked) begin // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 208:20]
      if (2'h0 == set) begin // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 210:18]
        if (2'h0 == step) begin // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 212:23]
          if (io_mixPc) begin // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 214:29]
            matrix_c_2 <= _matrix_c_2_T; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 218:29]
          end else begin
            matrix_c_2 <= _matrix_c_2_T_1; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 223:29]
          end
        end else if (2'h1 == step) begin // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 212:23]
          matrix_c_2 <= _GEN_3146;
        end else begin
          matrix_c_2 <= _GEN_3180;
        end
      end else if (2'h1 == set) begin // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 210:18]
        if (_T_1) begin // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 254:24]
          matrix_c_2 <= _GEN_3331;
        end else begin
          matrix_c_2 <= _GEN_3395;
        end
      end else if (2'h2 == set) begin // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 210:18]
        matrix_c_2 <= _GEN_3636;
      end else begin
        matrix_c_2 <= _GEN_3903;
      end
    end
    if (handshaked) begin // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 208:20]
      if (2'h0 == set) begin // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 210:18]
        if (2'h0 == step) begin // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 212:23]
          if (io_mixPc) begin // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 214:29]
            matrix_c_3 <= _matrix_c_3_T; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 218:29]
          end else begin
            matrix_c_3 <= _matrix_c_3_T_1; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 223:29]
          end
        end else if (2'h1 == step) begin // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 212:23]
          matrix_c_3 <= _GEN_4678;
        end else begin
          matrix_c_3 <= _GEN_4712;
        end
      end else if (2'h1 == set) begin // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 210:18]
        if (_T_1) begin // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 254:24]
          matrix_c_3 <= _GEN_4859;
        end else begin
          matrix_c_3 <= _GEN_4919;
        end
      end else if (2'h2 == set) begin // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 210:18]
        matrix_c_3 <= _GEN_5152;
      end else begin
        matrix_c_3 <= _GEN_5411;
      end
    end
    if (handshaked) begin // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 208:20]
      if (2'h0 == set) begin // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 210:18]
        if (2'h0 == step) begin // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 212:23]
          if (io_mixPc) begin // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 214:29]
            matrix_c_4 <= _matrix_c_4_T; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 218:29]
          end else begin
            matrix_c_4 <= _matrix_c_4_T_1; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 223:29]
          end
        end else if (2'h1 == step) begin // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 212:23]
          matrix_c_4 <= _GEN_6202;
        end else begin
          matrix_c_4 <= _GEN_6236;
        end
      end else if (2'h1 == set) begin // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 210:18]
        if (_T_1) begin // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 254:24]
          matrix_c_4 <= _GEN_6389;
        end else begin
          matrix_c_4 <= _GEN_6459;
        end
      end else if (2'h2 == set) begin // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 210:18]
        matrix_c_4 <= _GEN_6708;
      end else begin
        matrix_c_4 <= _GEN_6983;
      end
    end
    if (handshaked) begin // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 208:20]
      if (2'h0 == set) begin // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 210:18]
        if (2'h0 == step) begin // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 212:23]
          if (io_mixPc) begin // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 214:29]
            matrix_c_5 <= _matrix_c_5_T; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 218:29]
          end else begin
            matrix_c_5 <= _matrix_c_5_T_1; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 223:29]
          end
        end else if (2'h1 == step) begin // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 212:23]
          matrix_c_5 <= _GEN_7766;
        end else begin
          matrix_c_5 <= _GEN_7800;
        end
      end else if (2'h1 == set) begin // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 210:18]
        if (_T_1) begin // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 254:24]
          matrix_c_5 <= _GEN_7949;
        end else begin
          matrix_c_5 <= _GEN_8015;
        end
      end else if (2'h2 == set) begin // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 210:18]
        matrix_c_5 <= _GEN_8256;
      end else begin
        matrix_c_5 <= _GEN_8523;
      end
    end
    if (handshaked) begin // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 208:20]
      if (2'h0 == set) begin // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 210:18]
        if (2'h0 == step) begin // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 212:23]
          if (io_mixPc) begin // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 214:29]
            matrix_c_6 <= _matrix_c_6_T; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 218:29]
          end else begin
            matrix_c_6 <= _matrix_c_6_T_1; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 223:29]
          end
        end else if (2'h1 == step) begin // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 212:23]
          matrix_c_6 <= _GEN_9306;
        end else begin
          matrix_c_6 <= _GEN_9340;
        end
      end else if (2'h1 == set) begin // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 210:18]
        if (_T_1) begin // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 254:24]
          matrix_c_6 <= _GEN_9491;
        end else begin
          matrix_c_6 <= _GEN_9555;
        end
      end else if (2'h2 == set) begin // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 210:18]
        matrix_c_6 <= _GEN_9796;
      end else begin
        matrix_c_6 <= _GEN_10063;
      end
    end
    if (handshaked) begin // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 208:20]
      if (2'h0 == set) begin // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 210:18]
        if (2'h0 == step) begin // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 212:23]
          if (io_mixPc) begin // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 214:29]
            matrix_c_7 <= _matrix_c_7_T; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 218:29]
          end else begin
            matrix_c_7 <= _matrix_c_7_T_1; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 223:29]
          end
        end else if (2'h1 == step) begin // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 212:23]
          matrix_c_7 <= _GEN_10838;
        end else begin
          matrix_c_7 <= _GEN_10872;
        end
      end else if (2'h1 == set) begin // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 210:18]
        if (_T_1) begin // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 254:24]
          matrix_c_7 <= _GEN_11019;
        end else begin
          matrix_c_7 <= _GEN_11079;
        end
      end else if (2'h2 == set) begin // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 210:18]
        matrix_c_7 <= _GEN_11312;
      end else begin
        matrix_c_7 <= _GEN_11571;
      end
    end
    if (handshaked) begin // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 169:32]
      io_top_src_valid_r <= in_valid; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 169:32]
    end
    if (handshaked) begin // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 173:46]
      io_top_src_bits_ctrl_mixPcMode_r <= io_mixPc; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Manager.scala 173:46]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {2{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    rf[initvar] = _RAND_0[63:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  set = _RAND_1[1:0];
  _RAND_2 = {1{`RANDOM}};
  step = _RAND_2[1:0];
  _RAND_3 = {1{`RANDOM}};
  out_set = _RAND_3[1:0];
  _RAND_4 = {1{`RANDOM}};
  out_step = _RAND_4[1:0];
  _RAND_5 = {1{`RANDOM}};
  exec_en = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  tx_en = _RAND_6[0:0];
  _RAND_7 = {8{`RANDOM}};
  matrix_a_0 = _RAND_7[255:0];
  _RAND_8 = {8{`RANDOM}};
  matrix_a_1 = _RAND_8[255:0];
  _RAND_9 = {8{`RANDOM}};
  matrix_a_2 = _RAND_9[255:0];
  _RAND_10 = {8{`RANDOM}};
  matrix_a_3 = _RAND_10[255:0];
  _RAND_11 = {8{`RANDOM}};
  matrix_a_4 = _RAND_11[255:0];
  _RAND_12 = {8{`RANDOM}};
  matrix_a_5 = _RAND_12[255:0];
  _RAND_13 = {8{`RANDOM}};
  matrix_a_6 = _RAND_13[255:0];
  _RAND_14 = {8{`RANDOM}};
  matrix_a_7 = _RAND_14[255:0];
  _RAND_15 = {8{`RANDOM}};
  matrix_b_0 = _RAND_15[255:0];
  _RAND_16 = {8{`RANDOM}};
  matrix_b_1 = _RAND_16[255:0];
  _RAND_17 = {8{`RANDOM}};
  matrix_b_2 = _RAND_17[255:0];
  _RAND_18 = {8{`RANDOM}};
  matrix_b_3 = _RAND_18[255:0];
  _RAND_19 = {8{`RANDOM}};
  matrix_b_4 = _RAND_19[255:0];
  _RAND_20 = {8{`RANDOM}};
  matrix_b_5 = _RAND_20[255:0];
  _RAND_21 = {8{`RANDOM}};
  matrix_b_6 = _RAND_21[255:0];
  _RAND_22 = {8{`RANDOM}};
  matrix_b_7 = _RAND_22[255:0];
  _RAND_23 = {8{`RANDOM}};
  matrix_c_0 = _RAND_23[255:0];
  _RAND_24 = {8{`RANDOM}};
  matrix_c_1 = _RAND_24[255:0];
  _RAND_25 = {8{`RANDOM}};
  matrix_c_2 = _RAND_25[255:0];
  _RAND_26 = {8{`RANDOM}};
  matrix_c_3 = _RAND_26[255:0];
  _RAND_27 = {8{`RANDOM}};
  matrix_c_4 = _RAND_27[255:0];
  _RAND_28 = {8{`RANDOM}};
  matrix_c_5 = _RAND_28[255:0];
  _RAND_29 = {8{`RANDOM}};
  matrix_c_6 = _RAND_29[255:0];
  _RAND_30 = {8{`RANDOM}};
  matrix_c_7 = _RAND_30[255:0];
  _RAND_31 = {1{`RANDOM}};
  io_top_src_valid_r = _RAND_31[0:0];
  _RAND_32 = {1{`RANDOM}};
  io_top_src_bits_ctrl_mixPcMode_r = _RAND_32[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module LZC(
  input  [10:0] io_in, // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/LZC.scala 11:14]
  output [3:0]  io_out // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/LZC.scala 11:14]
);
  wire [3:0] _io_out_T_11 = io_in[1] ? 4'h9 : 4'ha; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [3:0] _io_out_T_12 = io_in[2] ? 4'h8 : _io_out_T_11; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [3:0] _io_out_T_13 = io_in[3] ? 4'h7 : _io_out_T_12; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [3:0] _io_out_T_14 = io_in[4] ? 4'h6 : _io_out_T_13; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [3:0] _io_out_T_15 = io_in[5] ? 4'h5 : _io_out_T_14; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [3:0] _io_out_T_16 = io_in[6] ? 4'h4 : _io_out_T_15; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [3:0] _io_out_T_17 = io_in[7] ? 4'h3 : _io_out_T_16; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [3:0] _io_out_T_18 = io_in[8] ? 4'h2 : _io_out_T_17; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [3:0] _io_out_T_19 = io_in[9] ? 4'h1 : _io_out_T_18; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  assign io_out = io_in[10] ? 4'h0 : _io_out_T_19; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
endmodule
module FMULnoRound(
  output        io_in_ready, // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FMUL.scala 26:14]
  input         io_in_valid, // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FMUL.scala 26:14]
  input  [15:0] io_in_bits_a, // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FMUL.scala 26:14]
  input  [15:0] io_in_bits_b, // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FMUL.scala 26:14]
  input         io_toFADD_ready, // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FMUL.scala 26:14]
  output        io_toFADD_valid, // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FMUL.scala 26:14]
  output [31:0] io_toFADD_bits_fp_prod, // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FMUL.scala 26:14]
  output        io_toFADD_bits_inter_flags_isNaN, // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FMUL.scala 26:14]
  output        io_toFADD_bits_inter_flags_isInf // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FMUL.scala 26:14]
);
  wire [10:0] aLZC_lzc_io_in; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/LZC.scala 21:21]
  wire [3:0] aLZC_lzc_io_out; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/LZC.scala 21:21]
  wire [10:0] bLZC_lzc_io_in; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/LZC.scala 21:21]
  wire [3:0] bLZC_lzc_io_out; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/LZC.scala 21:21]
  wire  fp_a_sign = io_in_bits_a[15]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/package.scala 58:19]
  wire [4:0] fp_a_exp = io_in_bits_a[14:10]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/package.scala 59:18]
  wire [9:0] fp_a_sig = io_in_bits_a[9:0]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/package.scala 60:18]
  wire  fp_b_sign = io_in_bits_b[15]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/package.scala 58:19]
  wire [4:0] fp_b_exp = io_in_bits_b[14:10]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/package.scala 59:18]
  wire [9:0] fp_b_sig = io_in_bits_b[9:0]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/package.scala 60:18]
  wire  expNotZero = |fp_a_exp; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/package.scala 31:28]
  wire  expIsOnes = &fp_a_exp; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/package.scala 32:27]
  wire  sigNotZero = |fp_a_sig; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/package.scala 33:28]
  wire  decode_a_expIsZero = ~expNotZero; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/package.scala 36:27]
  wire  decode_a_sigIsZero = ~sigNotZero; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/package.scala 39:27]
  wire  decode_a_isInf = expIsOnes & decode_a_sigIsZero; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/package.scala 41:40]
  wire  decode_a_isZero = decode_a_expIsZero & decode_a_sigIsZero; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/package.scala 42:41]
  wire  decode_a_isNaN = expIsOnes & sigNotZero; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/package.scala 43:40]
  wire  expNotZero_1 = |fp_b_exp; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/package.scala 31:28]
  wire  expIsOnes_1 = &fp_b_exp; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/package.scala 32:27]
  wire  sigNotZero_1 = |fp_b_sig; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/package.scala 33:28]
  wire  decode_b_expIsZero = ~expNotZero_1; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/package.scala 36:27]
  wire  decode_b_sigIsZero = ~sigNotZero_1; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/package.scala 39:27]
  wire  decode_b_isInf = expIsOnes_1 & decode_b_sigIsZero; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/package.scala 41:40]
  wire  decode_b_isZero = decode_b_expIsZero & decode_b_sigIsZero; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/package.scala 42:41]
  wire  decode_b_isNaN = expIsOnes_1 & sigNotZero_1; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/package.scala 43:40]
  wire  raw_a_isSub = sigNotZero & decode_a_expIsZero; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/package.scala 81:78]
  wire [4:0] _raw_a_inner_exp_T_1 = fp_a_exp + 5'h1; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/package.scala 83:38]
  wire [4:0] raw_a_exp = raw_a_isSub ? _raw_a_inner_exp_T_1 : fp_a_exp; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/package.scala 83:23]
  wire [10:0] raw_a_sig = {expNotZero,fp_a_sig}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/package.scala 84:23]
  wire  raw_b_isSub = sigNotZero_1 & decode_b_expIsZero; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/package.scala 81:78]
  wire [4:0] _raw_b_inner_exp_T_1 = fp_b_exp + 5'h1; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/package.scala 83:38]
  wire [4:0] raw_b_exp = raw_b_isSub ? _raw_b_inner_exp_T_1 : fp_b_exp; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/package.scala 83:23]
  wire [10:0] raw_b_sig = {expNotZero_1,fp_b_sig}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/package.scala 84:23]
  wire  hasZero = decode_a_isZero | decode_b_isZero; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FMUL.scala 39:33]
  wire  resultSign = fp_a_sign ^ fp_b_sign; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FMUL.scala 40:30]
  wire [5:0] _expSum_T = {1'h0,raw_a_exp}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FMUL.scala 41:19]
  wire [5:0] _expSum_T_1 = {1'h0,raw_b_exp}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FMUL.scala 41:46]
  wire [5:0] expSum = _expSum_T + _expSum_T_1; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FMUL.scala 41:41]
  wire [7:0] _expSumUpPc_T = {2'h0,expSum}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FMUL.scala 44:23]
  wire [7:0] expSumUpPc = _expSumUpPc_T + 8'h61; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FMUL.scala 44:71]
  wire [7:0] resultExpNoShift = hasZero ? 8'h0 : expSumUpPc; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [21:0] resultSigNoShift = raw_a_sig * raw_b_sig; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FMUL.scala 51:37]
  wire [3:0] lzcRaw = aLZC_lzc_io_out + bLZC_lzc_io_out; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FMUL.scala 57:21]
  wire [21:0] ErrorDetectMask = 22'h200000 >> lzcRaw; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FMUL.scala 58:68]
  wire [21:0] _lzcError_T = resultSigNoShift & ErrorDetectMask; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FMUL.scala 59:37]
  wire  lzcError = ~(|_lzcError_T); // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FMUL.scala 59:18]
  wire [3:0] _lzc_T_1 = lzcRaw + 4'h1; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FMUL.scala 60:34]
  wire [3:0] lzc = lzcError ? _lzc_T_1 : lzcRaw; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FMUL.scala 60:16]
  wire [7:0] _shiftLimit_T_1 = resultExpNoShift + 8'h1; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FMUL.scala 61:38]
  wire [7:0] _GEN_0 = {{4'd0}, lzc}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FMUL.scala 61:45]
  wire  shiftLimit = _shiftLimit_T_1 <= _GEN_0; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FMUL.scala 61:45]
  wire [7:0] _resultSigShifted_T = shiftLimit ? resultExpNoShift : {{4'd0}, lzc}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FMUL.scala 63:50]
  wire [276:0] _GEN_1 = {{255'd0}, resultSigNoShift}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FMUL.scala 63:44]
  wire [276:0] _resultSigShifted_T_1 = _GEN_1 << _resultSigShifted_T; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FMUL.scala 63:44]
  wire [21:0] resultSigShifted = _resultSigShifted_T_1[21:0]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FMUL.scala 63:86]
  wire [7:0] _resultExpShifted_T_1 = resultExpNoShift - _GEN_0; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FMUL.scala 64:79]
  wire [7:0] _resultExpShifted_T_3 = _resultExpShifted_T_1 + 8'h1; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FMUL.scala 64:85]
  wire [7:0] resultExpShifted = shiftLimit ? 8'h0 : _resultExpShifted_T_3; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FMUL.scala 64:29]
  wire  hasNaN = decode_a_isNaN | decode_b_isNaN; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FMUL.scala 68:31]
  wire  hasInf = decode_a_isInf | decode_b_isInf; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FMUL.scala 70:31]
  wire  special_case_happen = hasZero | hasNaN | hasInf; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FMUL.scala 71:47]
  wire  zero_mul_inf = hasZero & hasInf; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FMUL.scala 73:30]
  wire  nan_result = hasNaN | zero_mul_inf; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FMUL.scala 74:27]
  wire [31:0] _special_result_T_2 = {resultSign,8'hff,23'h0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FMUL.scala 79:10]
  wire [31:0] _special_result_T_3 = {resultSign,31'h0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FMUL.scala 83:10]
  wire [31:0] _special_result_T_4 = hasInf ? _special_result_T_2 : _special_result_T_3; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FMUL.scala 78:8]
  wire [31:0] special_result = nan_result ? 32'h7fc00000 : _special_result_T_4; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FMUL.scala 76:27]
  wire [31:0] _io_toFADD_bits_fp_prod_T_1 = {resultSign,resultExpShifted,resultSigShifted[20:0],2'h0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FMUL.scala 91:8]
  LZC aLZC_lzc ( // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/LZC.scala 21:21]
    .io_in(aLZC_lzc_io_in),
    .io_out(aLZC_lzc_io_out)
  );
  LZC bLZC_lzc ( // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/LZC.scala 21:21]
    .io_in(bLZC_lzc_io_in),
    .io_out(bLZC_lzc_io_out)
  );
  assign io_in_ready = io_toFADD_ready; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FMUL.scala 93:15]
  assign io_toFADD_valid = io_in_valid; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FMUL.scala 94:19]
  assign io_toFADD_bits_fp_prod = special_case_happen ? special_result : _io_toFADD_bits_fp_prod_T_1; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FMUL.scala 89:32]
  assign io_toFADD_bits_inter_flags_isNaN = hasNaN | zero_mul_inf; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FMUL.scala 74:27]
  assign io_toFADD_bits_inter_flags_isInf = decode_a_isInf | decode_b_isInf; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FMUL.scala 70:31]
  assign aLZC_lzc_io_in = {expNotZero,fp_a_sig}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/package.scala 84:23]
  assign bLZC_lzc_io_in = {expNotZero_1,fp_b_sig}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/package.scala 84:23]
endmodule
module LZC_8(
  input  [9:0] io_in, // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/LZC.scala 11:14]
  output [3:0] io_out // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/LZC.scala 11:14]
);
  wire [3:0] _io_out_T_10 = io_in[1] ? 4'h8 : 4'h9; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [3:0] _io_out_T_11 = io_in[2] ? 4'h7 : _io_out_T_10; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [3:0] _io_out_T_12 = io_in[3] ? 4'h6 : _io_out_T_11; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [3:0] _io_out_T_13 = io_in[4] ? 4'h5 : _io_out_T_12; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [3:0] _io_out_T_14 = io_in[5] ? 4'h4 : _io_out_T_13; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [3:0] _io_out_T_15 = io_in[6] ? 4'h3 : _io_out_T_14; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [3:0] _io_out_T_16 = io_in[7] ? 4'h2 : _io_out_T_15; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [3:0] _io_out_T_17 = io_in[8] ? 4'h1 : _io_out_T_16; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  assign io_out = io_in[9] ? 4'h0 : _io_out_T_17; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
endmodule
module FPUpConverter(
  output        io_in_ready, // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FPToFP.scala 246:14]
  input  [15:0] io_in_bits_in, // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FPToFP.scala 246:14]
  input         io_out_ready, // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FPToFP.scala 246:14]
  output [31:0] io_out_bits_result // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FPToFP.scala 246:14]
);
  wire [9:0] subnormal_shamt_lzc_io_in; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/LZC.scala 21:21]
  wire [3:0] subnormal_shamt_lzc_io_out; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/LZC.scala 21:21]
  wire  fp_in_sign = io_in_bits_in[15]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/package.scala 58:19]
  wire [4:0] fp_in_exp = io_in_bits_in[14:10]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/package.scala 59:18]
  wire [9:0] fp_in_sig = io_in_bits_in[9:0]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/package.scala 60:18]
  wire  decode_in_expNotZero = |fp_in_exp; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/package.scala 31:28]
  wire  decode_in_expIsOnes = &fp_in_exp; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/package.scala 32:27]
  wire  decode_in_sigNotZero = |fp_in_sig; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/package.scala 33:28]
  wire  decode_in__expIsZero = ~decode_in_expNotZero; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/package.scala 36:27]
  wire  decode_in__isSubnormal = decode_in__expIsZero & decode_in_sigNotZero; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/package.scala 40:46]
  wire  decode_in__isNaN = decode_in_expIsOnes & decode_in_sigNotZero; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/package.scala 43:40]
  wire [7:0] _GEN_0 = {{3'd0}, fp_in_exp}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FPToFP.scala 258:45]
  wire [7:0] normal_exp = 8'h70 + _GEN_0; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FPToFP.scala 258:45]
  wire [24:0] _GEN_2 = {{15'd0}, fp_in_sig}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FPToFP.scala 264:20]
  wire [24:0] _subnormal_sig_T = _GEN_2 << subnormal_shamt_lzc_io_out; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FPToFP.scala 264:20]
  wire [7:0] _GEN_1 = {{4'd0}, subnormal_shamt_lzc_io_out}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FPToFP.scala 265:48]
  wire [7:0] subnormal_exp = 8'h70 - _GEN_1; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FPToFP.scala 265:48]
  wire  _result_T_1 = ~decode_in__isNaN & fp_in_sign; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FPToFP.scala 270:22]
  wire  _result_T_4 = ~decode_in_expIsOnes & ~decode_in__expIsZero; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FPToFP.scala 276:30]
  wire [7:0] _result_T_6 = decode_in_expIsOnes ? 8'hff : 8'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [7:0] _result_T_8 = decode_in__isSubnormal ? subnormal_exp : 8'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [7:0] _result_T_9 = _result_T_4 ? normal_exp : 8'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [7:0] _result_T_11 = _result_T_6 | _result_T_8; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [7:0] _result_T_12 = _result_T_11 | _result_T_9; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [22:0] _result_T_16 = {decode_in_sigNotZero,22'h0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FPToFP.scala 292:12]
  wire [22:0] _result_T_17 = {_subnormal_sig_T[8:0],1'h0,13'h0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FPToFP.scala 293:12]
  wire [22:0] _result_T_18 = {fp_in_sig,13'h0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FPToFP.scala 294:12]
  wire [22:0] _result_T_19 = decode_in_expIsOnes ? _result_T_16 : 23'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [22:0] _result_T_20 = decode_in__expIsZero ? _result_T_17 : 23'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [22:0] _result_T_21 = _result_T_4 ? _result_T_18 : 23'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [22:0] _result_T_22 = _result_T_19 | _result_T_20; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [22:0] _result_T_23 = _result_T_22 | _result_T_21; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [8:0] result_hi = {_result_T_1,_result_T_12}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FPToFP.scala 269:19]
  LZC_8 subnormal_shamt_lzc ( // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/LZC.scala 21:21]
    .io_in(subnormal_shamt_lzc_io_in),
    .io_out(subnormal_shamt_lzc_io_out)
  );
  assign io_in_ready = io_out_ready; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FPToFP.scala 301:15]
  assign io_out_bits_result = {result_hi,_result_T_23}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FPToFP.scala 269:19]
  assign subnormal_shamt_lzc_io_in = io_in_bits_in[9:0]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/package.scala 60:18]
endmodule
module ShiftRightJam(
  input  [25:0] io_in, // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/ShiftRightJam.scala 11:14]
  input  [4:0]  io_shamt, // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/ShiftRightJam.scala 11:14]
  output [25:0] io_out, // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/ShiftRightJam.scala 11:14]
  output        io_sticky // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/ShiftRightJam.scala 11:14]
);
  wire  exceed_max_shift = io_shamt > 5'h1a; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/ShiftRightJam.scala 17:35]
  wire [31:0] _sticky_mask_T = 32'h1 << io_shamt; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/ShiftRightJam.scala 20:11]
  wire [31:0] _sticky_mask_T_2 = _sticky_mask_T - 32'h1; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/ShiftRightJam.scala 20:28]
  wire [25:0] _sticky_mask_T_5 = exceed_max_shift ? 26'h3ffffff : 26'h0; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/ShiftRightJam.scala 20:53]
  wire [25:0] sticky_mask = _sticky_mask_T_2[25:0] | _sticky_mask_T_5; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/ShiftRightJam.scala 20:47]
  wire [25:0] _io_out_T = io_in >> io_shamt; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/ShiftRightJam.scala 21:46]
  wire [25:0] _io_sticky_T = io_in & sticky_mask; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/ShiftRightJam.scala 22:23]
  assign io_out = exceed_max_shift ? 26'h0 : _io_out_T; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/ShiftRightJam.scala 21:16]
  assign io_sticky = |_io_sticky_T; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/ShiftRightJam.scala 22:38]
endmodule
module RoundingUnit(
  input  [22:0] io_in, // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/RoundingUnit.scala 7:14]
  input         io_roundIn, // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/RoundingUnit.scala 7:14]
  input         io_stickyIn, // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/RoundingUnit.scala 7:14]
  output [22:0] io_out, // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/RoundingUnit.scala 7:14]
  output        io_cout // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/RoundingUnit.scala 7:14]
);
  wire  g = io_in[0]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/RoundingUnit.scala 19:25]
  wire  r_up = io_roundIn & io_stickyIn | io_roundIn & ~io_stickyIn & g; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/RoundingUnit.scala 25:24]
  wire [22:0] out_r_up = io_in + 23'h1; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/RoundingUnit.scala 32:24]
  assign io_out = r_up ? out_r_up : io_in; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/RoundingUnit.scala 33:16]
  assign io_cout = r_up & &io_in; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/RoundingUnit.scala 36:19]
endmodule
module TininessRounder(
  input  [26:0] io_in_sig // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/RoundingUnit.scala 60:14]
);
  wire [22:0] rounder_io_in; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/RoundingUnit.scala 44:25]
  wire  rounder_io_roundIn; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/RoundingUnit.scala 44:25]
  wire  rounder_io_stickyIn; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/RoundingUnit.scala 44:25]
  wire [22:0] rounder_io_out; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/RoundingUnit.scala 44:25]
  wire  rounder_io_cout; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/RoundingUnit.scala 44:25]
  RoundingUnit rounder ( // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/RoundingUnit.scala 44:25]
    .io_in(rounder_io_in),
    .io_roundIn(rounder_io_roundIn),
    .io_stickyIn(rounder_io_stickyIn),
    .io_out(rounder_io_out),
    .io_cout(rounder_io_cout)
  );
  assign rounder_io_in = io_in_sig[24:2]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/RoundingUnit.scala 45:33]
  assign rounder_io_roundIn = io_in_sig[1]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/RoundingUnit.scala 46:50]
  assign rounder_io_stickyIn = |io_in_sig[0]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/RoundingUnit.scala 47:51]
endmodule
module FarPath(
  input         io_in_a_sign, // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FADD.scala 9:14]
  input  [7:0]  io_in_a_exp, // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FADD.scala 9:14]
  input  [23:0] io_in_a_sig, // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FADD.scala 9:14]
  input  [7:0]  io_in_b_exp, // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FADD.scala 9:14]
  input  [23:0] io_in_b_sig, // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FADD.scala 9:14]
  input         io_in_addSig, // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FADD.scala 9:14]
  input         io_in_tinyAdd, // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FADD.scala 9:14]
  input  [4:0]  io_in_shiftNum, // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FADD.scala 9:14]
  output [31:0] io_out_result, // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FADD.scala 9:14]
  output        io_out_far_path_of // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FADD.scala 9:14]
);
  wire [25:0] shiftRightJam_io_in; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/ShiftRightJam.scala 27:31]
  wire [4:0] shiftRightJam_io_shamt; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/ShiftRightJam.scala 27:31]
  wire [25:0] shiftRightJam_io_out; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/ShiftRightJam.scala 27:31]
  wire  shiftRightJam_io_sticky; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/ShiftRightJam.scala 27:31]
  wire [26:0] far_path_tininess_rounder_io_in_sig; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FADD.scala 73:41]
  wire [22:0] far_path_rounder_io_in; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/RoundingUnit.scala 44:25]
  wire  far_path_rounder_io_roundIn; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/RoundingUnit.scala 44:25]
  wire  far_path_rounder_io_stickyIn; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/RoundingUnit.scala 44:25]
  wire [22:0] far_path_rounder_io_out; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/RoundingUnit.scala 44:25]
  wire  far_path_rounder_io_cout; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/RoundingUnit.scala 44:25]
  wire  aIsZero = ~(|io_in_a_exp); // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FADD.scala 26:17]
  wire  bIsZero = ~(|io_in_b_exp); // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FADD.scala 27:17]
  wire  bothZero = aIsZero & bIsZero; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FADD.scala 28:26]
  wire [27:0] pos_sigB = {1'h0,shiftRightJam_io_out,shiftRightJam_io_sticky}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FADD.scala 33:21]
  wire [26:0] _neg_sigB_T = {shiftRightJam_io_out,shiftRightJam_io_sticky}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FADD.scala 34:36]
  wire [26:0] _neg_sigB_T_1 = ~_neg_sigB_T; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FADD.scala 34:32]
  wire [26:0] _neg_sigB_T_3 = _neg_sigB_T_1 + 27'h1; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FADD.scala 34:63]
  wire [27:0] neg_sigB = {1'h1,_neg_sigB_T_3}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FADD.scala 34:21]
  wire [27:0] adder_in_sigB = io_in_addSig ? pos_sigB : neg_sigB; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FADD.scala 35:26]
  wire [27:0] adder_in_sigA = {1'h0,io_in_a_sig,3'h0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FADD.scala 36:26]
  wire [27:0] resultSigInNormalCase = adder_in_sigA + adder_in_sigB; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FADD.scala 37:45]
  wire [27:0] result_sig_raw = bIsZero ? adder_in_sigA : resultSigInNormalCase; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FADD.scala 39:27]
  wire  cout = result_sig_raw[27]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FADD.scala 41:33]
  wire  keep = result_sig_raw[26]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FADD.scala 42:41]
  wire  _resultSigNoRound_T = keep | io_in_tinyAdd; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FADD.scala 45:19]
  wire [26:0] _resultSigNoRound_T_4 = {result_sig_raw[27:2],|result_sig_raw[1:0]}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FADD.scala 47:44]
  wire [26:0] _resultSigNoRound_T_9 = {result_sig_raw[26:1],|result_sig_raw[0]}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FADD.scala 48:52]
  wire [26:0] _resultSigNoRound_T_14 = {result_sig_raw[25:0],1'h0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FADD.scala 49:52]
  wire [26:0] _resultSigNoRound_T_15 = _resultSigNoRound_T ? _resultSigNoRound_T_9 : _resultSigNoRound_T_14; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [26:0] resultSigNoRound = cout ? _resultSigNoRound_T_4 : _resultSigNoRound_T_15; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [7:0] _resultExpNoRound_T_1 = io_in_a_exp + 8'h1; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FADD.scala 55:28]
  wire  _resultExpNoRound_T_2 = keep | bothZero; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FADD.scala 56:13]
  wire [7:0] _resultExpNoRound_T_5 = io_in_a_exp - 8'h1; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FADD.scala 57:43]
  wire [7:0] _resultExpNoRound_T_6 = _resultExpNoRound_T_2 ? io_in_a_exp : _resultExpNoRound_T_5; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [7:0] resultExpNoRound = cout ? _resultExpNoRound_T_1 : _resultExpNoRound_T_6; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [7:0] _GEN_0 = {{7'd0}, far_path_rounder_io_cout}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FADD.scala 85:55]
  wire [7:0] far_path_exp_rounded = _GEN_0 + resultExpNoRound; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FADD.scala 85:55]
  wire  far_path_may_of = &io_in_b_exp & io_in_addSig; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FADD.scala 88:42]
  wire  far_path_of_before_round = resultExpNoRound == 8'hff; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FADD.scala 93:22]
  wire  _far_path_of_after_round_T = resultExpNoRound == 8'hfe; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FADD.scala 95:22]
  wire  far_path_of_after_round = far_path_rounder_io_cout & _far_path_of_after_round_T; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FADD.scala 94:58]
  wire [8:0] io_out_result_hi = {io_in_a_sign,far_path_exp_rounded}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FADD.scala 103:8]
  ShiftRightJam shiftRightJam ( // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/ShiftRightJam.scala 27:31]
    .io_in(shiftRightJam_io_in),
    .io_shamt(shiftRightJam_io_shamt),
    .io_out(shiftRightJam_io_out),
    .io_sticky(shiftRightJam_io_sticky)
  );
  TininessRounder far_path_tininess_rounder ( // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FADD.scala 73:41]
    .io_in_sig(far_path_tininess_rounder_io_in_sig)
  );
  RoundingUnit far_path_rounder ( // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/RoundingUnit.scala 44:25]
    .io_in(far_path_rounder_io_in),
    .io_roundIn(far_path_rounder_io_roundIn),
    .io_stickyIn(far_path_rounder_io_stickyIn),
    .io_out(far_path_rounder_io_out),
    .io_cout(far_path_rounder_io_cout)
  );
  assign io_out_result = {io_out_result_hi,far_path_rounder_io_out}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FADD.scala 103:8]
  assign io_out_far_path_of = far_path_of_before_round | far_path_of_after_round | far_path_may_of; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FADD.scala 98:57]
  assign shiftRightJam_io_in = {io_in_b_sig,2'h0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FADD.scala 30:53]
  assign shiftRightJam_io_shamt = io_in_shiftNum; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/ShiftRightJam.scala 29:28]
  assign far_path_tininess_rounder_io_in_sig = cout ? _resultSigNoRound_T_4 : _resultSigNoRound_T_15; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  assign far_path_rounder_io_in = resultSigNoRound[25:3]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/RoundingUnit.scala 45:33]
  assign far_path_rounder_io_roundIn = resultSigNoRound[2]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/RoundingUnit.scala 46:50]
  assign far_path_rounder_io_stickyIn = |resultSigNoRound[1:0]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/RoundingUnit.scala 47:51]
endmodule
module PreEncoder(
  input  [24:0] io_g, // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/PreEncoder.scala 11:14]
  input  [24:0] io_s, // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/PreEncoder.scala 11:14]
  input  [24:0] io_e, // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/PreEncoder.scala 11:14]
  output [24:0] io_f // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/PreEncoder.scala 11:14]
);
  wire  _f_0_T_6 = ~io_e[1] & io_s[0]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/PreEncoder.scala 17:25]
  wire  _f_0_T_7 = io_e[1] & io_g[0] | _f_0_T_6; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/PreEncoder.scala 16:33]
  wire  _f_0_T_10 = io_e[1] & io_s[0]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/PreEncoder.scala 18:25]
  wire  _f_0_T_11 = _f_0_T_7 | _f_0_T_10; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/PreEncoder.scala 17:33]
  wire  f_0 = _f_0_T_11 | io_e[1] & io_s[0]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/PreEncoder.scala 18:33]
  wire  _f_1_T_4 = ~io_s[0]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/PreEncoder.scala 23:33]
  wire  _f_1_T_7 = ~io_e[2]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/PreEncoder.scala 24:14]
  wire  _f_1_T_12 = ~io_e[2] & io_s[1] & _f_1_T_4; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/PreEncoder.scala 24:30]
  wire  _f_1_T_13 = io_e[2] & io_g[1] & ~io_s[0] | _f_1_T_12; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/PreEncoder.scala 23:43]
  wire  _f_1_T_18 = ~io_g[0]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/PreEncoder.scala 25:33]
  wire  _f_1_T_19 = io_e[2] & io_s[1] & ~io_g[0]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/PreEncoder.scala 25:30]
  wire  _f_1_T_20 = _f_1_T_13 | _f_1_T_19; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/PreEncoder.scala 24:43]
  wire  _f_1_T_27 = _f_1_T_7 & io_g[1] & _f_1_T_18; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/PreEncoder.scala 26:30]
  wire  f_1 = _f_1_T_20 | _f_1_T_27; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/PreEncoder.scala 25:43]
  wire  _f_2_T_4 = ~io_s[1]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/PreEncoder.scala 23:33]
  wire  _f_2_T_7 = ~io_e[3]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/PreEncoder.scala 24:14]
  wire  _f_2_T_12 = ~io_e[3] & io_s[2] & _f_2_T_4; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/PreEncoder.scala 24:30]
  wire  _f_2_T_13 = io_e[3] & io_g[2] & ~io_s[1] | _f_2_T_12; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/PreEncoder.scala 23:43]
  wire  _f_2_T_18 = ~io_g[1]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/PreEncoder.scala 25:33]
  wire  _f_2_T_19 = io_e[3] & io_s[2] & ~io_g[1]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/PreEncoder.scala 25:30]
  wire  _f_2_T_20 = _f_2_T_13 | _f_2_T_19; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/PreEncoder.scala 24:43]
  wire  _f_2_T_27 = _f_2_T_7 & io_g[2] & _f_2_T_18; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/PreEncoder.scala 26:30]
  wire  f_2 = _f_2_T_20 | _f_2_T_27; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/PreEncoder.scala 25:43]
  wire  _f_3_T_4 = ~io_s[2]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/PreEncoder.scala 23:33]
  wire  _f_3_T_7 = ~io_e[4]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/PreEncoder.scala 24:14]
  wire  _f_3_T_12 = ~io_e[4] & io_s[3] & _f_3_T_4; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/PreEncoder.scala 24:30]
  wire  _f_3_T_13 = io_e[4] & io_g[3] & ~io_s[2] | _f_3_T_12; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/PreEncoder.scala 23:43]
  wire  _f_3_T_18 = ~io_g[2]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/PreEncoder.scala 25:33]
  wire  _f_3_T_19 = io_e[4] & io_s[3] & ~io_g[2]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/PreEncoder.scala 25:30]
  wire  _f_3_T_20 = _f_3_T_13 | _f_3_T_19; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/PreEncoder.scala 24:43]
  wire  _f_3_T_27 = _f_3_T_7 & io_g[3] & _f_3_T_18; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/PreEncoder.scala 26:30]
  wire  f_3 = _f_3_T_20 | _f_3_T_27; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/PreEncoder.scala 25:43]
  wire  _f_4_T_4 = ~io_s[3]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/PreEncoder.scala 23:33]
  wire  _f_4_T_7 = ~io_e[5]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/PreEncoder.scala 24:14]
  wire  _f_4_T_12 = ~io_e[5] & io_s[4] & _f_4_T_4; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/PreEncoder.scala 24:30]
  wire  _f_4_T_13 = io_e[5] & io_g[4] & ~io_s[3] | _f_4_T_12; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/PreEncoder.scala 23:43]
  wire  _f_4_T_18 = ~io_g[3]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/PreEncoder.scala 25:33]
  wire  _f_4_T_19 = io_e[5] & io_s[4] & ~io_g[3]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/PreEncoder.scala 25:30]
  wire  _f_4_T_20 = _f_4_T_13 | _f_4_T_19; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/PreEncoder.scala 24:43]
  wire  _f_4_T_27 = _f_4_T_7 & io_g[4] & _f_4_T_18; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/PreEncoder.scala 26:30]
  wire  f_4 = _f_4_T_20 | _f_4_T_27; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/PreEncoder.scala 25:43]
  wire  _f_5_T_4 = ~io_s[4]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/PreEncoder.scala 23:33]
  wire  _f_5_T_7 = ~io_e[6]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/PreEncoder.scala 24:14]
  wire  _f_5_T_12 = ~io_e[6] & io_s[5] & _f_5_T_4; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/PreEncoder.scala 24:30]
  wire  _f_5_T_13 = io_e[6] & io_g[5] & ~io_s[4] | _f_5_T_12; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/PreEncoder.scala 23:43]
  wire  _f_5_T_18 = ~io_g[4]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/PreEncoder.scala 25:33]
  wire  _f_5_T_19 = io_e[6] & io_s[5] & ~io_g[4]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/PreEncoder.scala 25:30]
  wire  _f_5_T_20 = _f_5_T_13 | _f_5_T_19; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/PreEncoder.scala 24:43]
  wire  _f_5_T_27 = _f_5_T_7 & io_g[5] & _f_5_T_18; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/PreEncoder.scala 26:30]
  wire  f_5 = _f_5_T_20 | _f_5_T_27; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/PreEncoder.scala 25:43]
  wire  _f_6_T_4 = ~io_s[5]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/PreEncoder.scala 23:33]
  wire  _f_6_T_7 = ~io_e[7]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/PreEncoder.scala 24:14]
  wire  _f_6_T_12 = ~io_e[7] & io_s[6] & _f_6_T_4; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/PreEncoder.scala 24:30]
  wire  _f_6_T_13 = io_e[7] & io_g[6] & ~io_s[5] | _f_6_T_12; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/PreEncoder.scala 23:43]
  wire  _f_6_T_18 = ~io_g[5]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/PreEncoder.scala 25:33]
  wire  _f_6_T_19 = io_e[7] & io_s[6] & ~io_g[5]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/PreEncoder.scala 25:30]
  wire  _f_6_T_20 = _f_6_T_13 | _f_6_T_19; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/PreEncoder.scala 24:43]
  wire  _f_6_T_27 = _f_6_T_7 & io_g[6] & _f_6_T_18; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/PreEncoder.scala 26:30]
  wire  f_6 = _f_6_T_20 | _f_6_T_27; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/PreEncoder.scala 25:43]
  wire  _f_7_T_4 = ~io_s[6]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/PreEncoder.scala 23:33]
  wire  _f_7_T_7 = ~io_e[8]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/PreEncoder.scala 24:14]
  wire  _f_7_T_12 = ~io_e[8] & io_s[7] & _f_7_T_4; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/PreEncoder.scala 24:30]
  wire  _f_7_T_13 = io_e[8] & io_g[7] & ~io_s[6] | _f_7_T_12; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/PreEncoder.scala 23:43]
  wire  _f_7_T_18 = ~io_g[6]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/PreEncoder.scala 25:33]
  wire  _f_7_T_19 = io_e[8] & io_s[7] & ~io_g[6]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/PreEncoder.scala 25:30]
  wire  _f_7_T_20 = _f_7_T_13 | _f_7_T_19; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/PreEncoder.scala 24:43]
  wire  _f_7_T_27 = _f_7_T_7 & io_g[7] & _f_7_T_18; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/PreEncoder.scala 26:30]
  wire  f_7 = _f_7_T_20 | _f_7_T_27; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/PreEncoder.scala 25:43]
  wire  _f_8_T_4 = ~io_s[7]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/PreEncoder.scala 23:33]
  wire  _f_8_T_7 = ~io_e[9]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/PreEncoder.scala 24:14]
  wire  _f_8_T_12 = ~io_e[9] & io_s[8] & _f_8_T_4; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/PreEncoder.scala 24:30]
  wire  _f_8_T_13 = io_e[9] & io_g[8] & ~io_s[7] | _f_8_T_12; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/PreEncoder.scala 23:43]
  wire  _f_8_T_18 = ~io_g[7]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/PreEncoder.scala 25:33]
  wire  _f_8_T_19 = io_e[9] & io_s[8] & ~io_g[7]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/PreEncoder.scala 25:30]
  wire  _f_8_T_20 = _f_8_T_13 | _f_8_T_19; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/PreEncoder.scala 24:43]
  wire  _f_8_T_27 = _f_8_T_7 & io_g[8] & _f_8_T_18; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/PreEncoder.scala 26:30]
  wire  f_8 = _f_8_T_20 | _f_8_T_27; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/PreEncoder.scala 25:43]
  wire  _f_9_T_4 = ~io_s[8]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/PreEncoder.scala 23:33]
  wire  _f_9_T_7 = ~io_e[10]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/PreEncoder.scala 24:14]
  wire  _f_9_T_12 = ~io_e[10] & io_s[9] & _f_9_T_4; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/PreEncoder.scala 24:30]
  wire  _f_9_T_13 = io_e[10] & io_g[9] & ~io_s[8] | _f_9_T_12; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/PreEncoder.scala 23:43]
  wire  _f_9_T_18 = ~io_g[8]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/PreEncoder.scala 25:33]
  wire  _f_9_T_19 = io_e[10] & io_s[9] & ~io_g[8]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/PreEncoder.scala 25:30]
  wire  _f_9_T_20 = _f_9_T_13 | _f_9_T_19; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/PreEncoder.scala 24:43]
  wire  _f_9_T_27 = _f_9_T_7 & io_g[9] & _f_9_T_18; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/PreEncoder.scala 26:30]
  wire  f_9 = _f_9_T_20 | _f_9_T_27; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/PreEncoder.scala 25:43]
  wire  _f_10_T_4 = ~io_s[9]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/PreEncoder.scala 23:33]
  wire  _f_10_T_7 = ~io_e[11]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/PreEncoder.scala 24:14]
  wire  _f_10_T_12 = ~io_e[11] & io_s[10] & _f_10_T_4; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/PreEncoder.scala 24:30]
  wire  _f_10_T_13 = io_e[11] & io_g[10] & ~io_s[9] | _f_10_T_12; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/PreEncoder.scala 23:43]
  wire  _f_10_T_18 = ~io_g[9]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/PreEncoder.scala 25:33]
  wire  _f_10_T_19 = io_e[11] & io_s[10] & ~io_g[9]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/PreEncoder.scala 25:30]
  wire  _f_10_T_20 = _f_10_T_13 | _f_10_T_19; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/PreEncoder.scala 24:43]
  wire  _f_10_T_27 = _f_10_T_7 & io_g[10] & _f_10_T_18; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/PreEncoder.scala 26:30]
  wire  f_10 = _f_10_T_20 | _f_10_T_27; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/PreEncoder.scala 25:43]
  wire  _f_11_T_4 = ~io_s[10]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/PreEncoder.scala 23:33]
  wire  _f_11_T_7 = ~io_e[12]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/PreEncoder.scala 24:14]
  wire  _f_11_T_12 = ~io_e[12] & io_s[11] & _f_11_T_4; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/PreEncoder.scala 24:30]
  wire  _f_11_T_13 = io_e[12] & io_g[11] & ~io_s[10] | _f_11_T_12; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/PreEncoder.scala 23:43]
  wire  _f_11_T_18 = ~io_g[10]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/PreEncoder.scala 25:33]
  wire  _f_11_T_19 = io_e[12] & io_s[11] & ~io_g[10]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/PreEncoder.scala 25:30]
  wire  _f_11_T_20 = _f_11_T_13 | _f_11_T_19; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/PreEncoder.scala 24:43]
  wire  _f_11_T_27 = _f_11_T_7 & io_g[11] & _f_11_T_18; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/PreEncoder.scala 26:30]
  wire  f_11 = _f_11_T_20 | _f_11_T_27; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/PreEncoder.scala 25:43]
  wire  _f_12_T_4 = ~io_s[11]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/PreEncoder.scala 23:33]
  wire  _f_12_T_7 = ~io_e[13]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/PreEncoder.scala 24:14]
  wire  _f_12_T_12 = ~io_e[13] & io_s[12] & _f_12_T_4; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/PreEncoder.scala 24:30]
  wire  _f_12_T_13 = io_e[13] & io_g[12] & ~io_s[11] | _f_12_T_12; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/PreEncoder.scala 23:43]
  wire  _f_12_T_18 = ~io_g[11]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/PreEncoder.scala 25:33]
  wire  _f_12_T_19 = io_e[13] & io_s[12] & ~io_g[11]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/PreEncoder.scala 25:30]
  wire  _f_12_T_20 = _f_12_T_13 | _f_12_T_19; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/PreEncoder.scala 24:43]
  wire  _f_12_T_27 = _f_12_T_7 & io_g[12] & _f_12_T_18; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/PreEncoder.scala 26:30]
  wire  f_12 = _f_12_T_20 | _f_12_T_27; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/PreEncoder.scala 25:43]
  wire  _f_13_T_4 = ~io_s[12]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/PreEncoder.scala 23:33]
  wire  _f_13_T_7 = ~io_e[14]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/PreEncoder.scala 24:14]
  wire  _f_13_T_12 = ~io_e[14] & io_s[13] & _f_13_T_4; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/PreEncoder.scala 24:30]
  wire  _f_13_T_13 = io_e[14] & io_g[13] & ~io_s[12] | _f_13_T_12; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/PreEncoder.scala 23:43]
  wire  _f_13_T_18 = ~io_g[12]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/PreEncoder.scala 25:33]
  wire  _f_13_T_19 = io_e[14] & io_s[13] & ~io_g[12]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/PreEncoder.scala 25:30]
  wire  _f_13_T_20 = _f_13_T_13 | _f_13_T_19; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/PreEncoder.scala 24:43]
  wire  _f_13_T_27 = _f_13_T_7 & io_g[13] & _f_13_T_18; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/PreEncoder.scala 26:30]
  wire  f_13 = _f_13_T_20 | _f_13_T_27; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/PreEncoder.scala 25:43]
  wire  _f_14_T_4 = ~io_s[13]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/PreEncoder.scala 23:33]
  wire  _f_14_T_7 = ~io_e[15]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/PreEncoder.scala 24:14]
  wire  _f_14_T_12 = ~io_e[15] & io_s[14] & _f_14_T_4; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/PreEncoder.scala 24:30]
  wire  _f_14_T_13 = io_e[15] & io_g[14] & ~io_s[13] | _f_14_T_12; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/PreEncoder.scala 23:43]
  wire  _f_14_T_18 = ~io_g[13]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/PreEncoder.scala 25:33]
  wire  _f_14_T_19 = io_e[15] & io_s[14] & ~io_g[13]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/PreEncoder.scala 25:30]
  wire  _f_14_T_20 = _f_14_T_13 | _f_14_T_19; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/PreEncoder.scala 24:43]
  wire  _f_14_T_27 = _f_14_T_7 & io_g[14] & _f_14_T_18; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/PreEncoder.scala 26:30]
  wire  f_14 = _f_14_T_20 | _f_14_T_27; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/PreEncoder.scala 25:43]
  wire  _f_15_T_4 = ~io_s[14]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/PreEncoder.scala 23:33]
  wire  _f_15_T_7 = ~io_e[16]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/PreEncoder.scala 24:14]
  wire  _f_15_T_12 = ~io_e[16] & io_s[15] & _f_15_T_4; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/PreEncoder.scala 24:30]
  wire  _f_15_T_13 = io_e[16] & io_g[15] & ~io_s[14] | _f_15_T_12; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/PreEncoder.scala 23:43]
  wire  _f_15_T_18 = ~io_g[14]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/PreEncoder.scala 25:33]
  wire  _f_15_T_19 = io_e[16] & io_s[15] & ~io_g[14]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/PreEncoder.scala 25:30]
  wire  _f_15_T_20 = _f_15_T_13 | _f_15_T_19; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/PreEncoder.scala 24:43]
  wire  _f_15_T_27 = _f_15_T_7 & io_g[15] & _f_15_T_18; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/PreEncoder.scala 26:30]
  wire  f_15 = _f_15_T_20 | _f_15_T_27; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/PreEncoder.scala 25:43]
  wire  _f_16_T_4 = ~io_s[15]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/PreEncoder.scala 23:33]
  wire  _f_16_T_7 = ~io_e[17]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/PreEncoder.scala 24:14]
  wire  _f_16_T_12 = ~io_e[17] & io_s[16] & _f_16_T_4; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/PreEncoder.scala 24:30]
  wire  _f_16_T_13 = io_e[17] & io_g[16] & ~io_s[15] | _f_16_T_12; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/PreEncoder.scala 23:43]
  wire  _f_16_T_18 = ~io_g[15]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/PreEncoder.scala 25:33]
  wire  _f_16_T_19 = io_e[17] & io_s[16] & ~io_g[15]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/PreEncoder.scala 25:30]
  wire  _f_16_T_20 = _f_16_T_13 | _f_16_T_19; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/PreEncoder.scala 24:43]
  wire  _f_16_T_27 = _f_16_T_7 & io_g[16] & _f_16_T_18; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/PreEncoder.scala 26:30]
  wire  f_16 = _f_16_T_20 | _f_16_T_27; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/PreEncoder.scala 25:43]
  wire  _f_17_T_4 = ~io_s[16]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/PreEncoder.scala 23:33]
  wire  _f_17_T_7 = ~io_e[18]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/PreEncoder.scala 24:14]
  wire  _f_17_T_12 = ~io_e[18] & io_s[17] & _f_17_T_4; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/PreEncoder.scala 24:30]
  wire  _f_17_T_13 = io_e[18] & io_g[17] & ~io_s[16] | _f_17_T_12; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/PreEncoder.scala 23:43]
  wire  _f_17_T_18 = ~io_g[16]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/PreEncoder.scala 25:33]
  wire  _f_17_T_19 = io_e[18] & io_s[17] & ~io_g[16]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/PreEncoder.scala 25:30]
  wire  _f_17_T_20 = _f_17_T_13 | _f_17_T_19; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/PreEncoder.scala 24:43]
  wire  _f_17_T_27 = _f_17_T_7 & io_g[17] & _f_17_T_18; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/PreEncoder.scala 26:30]
  wire  f_17 = _f_17_T_20 | _f_17_T_27; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/PreEncoder.scala 25:43]
  wire  _f_18_T_4 = ~io_s[17]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/PreEncoder.scala 23:33]
  wire  _f_18_T_7 = ~io_e[19]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/PreEncoder.scala 24:14]
  wire  _f_18_T_12 = ~io_e[19] & io_s[18] & _f_18_T_4; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/PreEncoder.scala 24:30]
  wire  _f_18_T_13 = io_e[19] & io_g[18] & ~io_s[17] | _f_18_T_12; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/PreEncoder.scala 23:43]
  wire  _f_18_T_18 = ~io_g[17]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/PreEncoder.scala 25:33]
  wire  _f_18_T_19 = io_e[19] & io_s[18] & ~io_g[17]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/PreEncoder.scala 25:30]
  wire  _f_18_T_20 = _f_18_T_13 | _f_18_T_19; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/PreEncoder.scala 24:43]
  wire  _f_18_T_27 = _f_18_T_7 & io_g[18] & _f_18_T_18; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/PreEncoder.scala 26:30]
  wire  f_18 = _f_18_T_20 | _f_18_T_27; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/PreEncoder.scala 25:43]
  wire  _f_19_T_4 = ~io_s[18]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/PreEncoder.scala 23:33]
  wire  _f_19_T_7 = ~io_e[20]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/PreEncoder.scala 24:14]
  wire  _f_19_T_12 = ~io_e[20] & io_s[19] & _f_19_T_4; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/PreEncoder.scala 24:30]
  wire  _f_19_T_13 = io_e[20] & io_g[19] & ~io_s[18] | _f_19_T_12; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/PreEncoder.scala 23:43]
  wire  _f_19_T_18 = ~io_g[18]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/PreEncoder.scala 25:33]
  wire  _f_19_T_19 = io_e[20] & io_s[19] & ~io_g[18]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/PreEncoder.scala 25:30]
  wire  _f_19_T_20 = _f_19_T_13 | _f_19_T_19; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/PreEncoder.scala 24:43]
  wire  _f_19_T_27 = _f_19_T_7 & io_g[19] & _f_19_T_18; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/PreEncoder.scala 26:30]
  wire  f_19 = _f_19_T_20 | _f_19_T_27; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/PreEncoder.scala 25:43]
  wire  _f_20_T_4 = ~io_s[19]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/PreEncoder.scala 23:33]
  wire  _f_20_T_7 = ~io_e[21]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/PreEncoder.scala 24:14]
  wire  _f_20_T_12 = ~io_e[21] & io_s[20] & _f_20_T_4; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/PreEncoder.scala 24:30]
  wire  _f_20_T_13 = io_e[21] & io_g[20] & ~io_s[19] | _f_20_T_12; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/PreEncoder.scala 23:43]
  wire  _f_20_T_18 = ~io_g[19]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/PreEncoder.scala 25:33]
  wire  _f_20_T_19 = io_e[21] & io_s[20] & ~io_g[19]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/PreEncoder.scala 25:30]
  wire  _f_20_T_20 = _f_20_T_13 | _f_20_T_19; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/PreEncoder.scala 24:43]
  wire  _f_20_T_27 = _f_20_T_7 & io_g[20] & _f_20_T_18; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/PreEncoder.scala 26:30]
  wire  f_20 = _f_20_T_20 | _f_20_T_27; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/PreEncoder.scala 25:43]
  wire  _f_21_T_4 = ~io_s[20]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/PreEncoder.scala 23:33]
  wire  _f_21_T_7 = ~io_e[22]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/PreEncoder.scala 24:14]
  wire  _f_21_T_12 = ~io_e[22] & io_s[21] & _f_21_T_4; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/PreEncoder.scala 24:30]
  wire  _f_21_T_13 = io_e[22] & io_g[21] & ~io_s[20] | _f_21_T_12; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/PreEncoder.scala 23:43]
  wire  _f_21_T_18 = ~io_g[20]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/PreEncoder.scala 25:33]
  wire  _f_21_T_19 = io_e[22] & io_s[21] & ~io_g[20]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/PreEncoder.scala 25:30]
  wire  _f_21_T_20 = _f_21_T_13 | _f_21_T_19; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/PreEncoder.scala 24:43]
  wire  _f_21_T_27 = _f_21_T_7 & io_g[21] & _f_21_T_18; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/PreEncoder.scala 26:30]
  wire  f_21 = _f_21_T_20 | _f_21_T_27; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/PreEncoder.scala 25:43]
  wire  _f_22_T_4 = ~io_s[21]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/PreEncoder.scala 23:33]
  wire  _f_22_T_7 = ~io_e[23]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/PreEncoder.scala 24:14]
  wire  _f_22_T_12 = ~io_e[23] & io_s[22] & _f_22_T_4; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/PreEncoder.scala 24:30]
  wire  _f_22_T_13 = io_e[23] & io_g[22] & ~io_s[21] | _f_22_T_12; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/PreEncoder.scala 23:43]
  wire  _f_22_T_18 = ~io_g[21]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/PreEncoder.scala 25:33]
  wire  _f_22_T_19 = io_e[23] & io_s[22] & ~io_g[21]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/PreEncoder.scala 25:30]
  wire  _f_22_T_20 = _f_22_T_13 | _f_22_T_19; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/PreEncoder.scala 24:43]
  wire  _f_22_T_27 = _f_22_T_7 & io_g[22] & _f_22_T_18; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/PreEncoder.scala 26:30]
  wire  f_22 = _f_22_T_20 | _f_22_T_27; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/PreEncoder.scala 25:43]
  wire  _f_23_T_4 = ~io_s[22]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/PreEncoder.scala 23:33]
  wire  _f_23_T_7 = ~io_e[24]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/PreEncoder.scala 24:14]
  wire  _f_23_T_12 = ~io_e[24] & io_s[23] & _f_23_T_4; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/PreEncoder.scala 24:30]
  wire  _f_23_T_13 = io_e[24] & io_g[23] & ~io_s[22] | _f_23_T_12; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/PreEncoder.scala 23:43]
  wire  _f_23_T_18 = ~io_g[22]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/PreEncoder.scala 25:33]
  wire  _f_23_T_19 = io_e[24] & io_s[23] & ~io_g[22]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/PreEncoder.scala 25:30]
  wire  _f_23_T_20 = _f_23_T_13 | _f_23_T_19; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/PreEncoder.scala 24:43]
  wire  _f_23_T_27 = _f_23_T_7 & io_g[23] & _f_23_T_18; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/PreEncoder.scala 26:30]
  wire  f_23 = _f_23_T_20 | _f_23_T_27; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/PreEncoder.scala 25:43]
  wire  f_24 = io_g[24] & ~io_s[23] | io_s[24] & ~io_g[23]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/PreEncoder.scala 21:36]
  wire [5:0] io_f_lo_lo = {f_5,f_4,f_3,f_2,f_1,f_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/PreEncoder.scala 29:14]
  wire [11:0] io_f_lo = {f_11,f_10,f_9,f_8,f_7,f_6,io_f_lo_lo}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/PreEncoder.scala 29:14]
  wire [5:0] io_f_hi_lo = {f_17,f_16,f_15,f_14,f_13,f_12}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/PreEncoder.scala 29:14]
  wire [12:0] io_f_hi = {f_24,f_23,f_22,f_21,f_20,f_19,f_18,io_f_hi_lo}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/PreEncoder.scala 29:14]
  assign io_f = {io_f_hi,io_f_lo}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/PreEncoder.scala 29:14]
endmodule
module node(
  input  [2:0] io_in_0, // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/node.scala 7:14]
  input  [2:0] io_in_2, // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/node.scala 7:14]
  output [1:0] io_out_0, // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/node.scala 7:14]
  output [1:0] io_out_2 // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/node.scala 7:14]
);
  wire  pout_0 = io_in_0[0] | io_in_2[0] & io_in_0[1]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/node.scala 16:19]
  wire  _pout_1_T_7 = io_in_2[0] | io_in_2[1]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/node.scala 17:47]
  wire  pout_1 = ~io_in_2[0] & io_in_0[1] | io_in_0[2] & (io_in_2[0] | io_in_2[1]); // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/node.scala 17:31]
  wire  zout_0 = io_in_2[0] & io_in_2[1]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/node.scala 18:19]
  wire  zout_1 = io_in_2[2] & _pout_1_T_7; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/node.scala 19:19]
  assign io_out_0 = {pout_1,pout_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/node.scala 22:19]
  assign io_out_2 = {zout_1,zout_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/node.scala 24:19]
endmodule
module ErrorDetector(
  input  [24:0] io_g, // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 12:14]
  input  [24:0] io_s, // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 12:14]
  input  [24:0] io_e, // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 12:14]
  output        io_y // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 12:14]
);
  wire [2:0] y_node0_io_in_0; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 31:23]
  wire [2:0] y_node0_io_in_2; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 31:23]
  wire [1:0] y_node0_io_out_0; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 31:23]
  wire [1:0] y_node0_io_out_2; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 31:23]
  wire [2:0] y_node_io_in_0; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 40:26]
  wire [2:0] y_node_io_in_2; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 40:26]
  wire [1:0] y_node_io_out_0; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 40:26]
  wire [1:0] y_node_io_out_2; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 40:26]
  wire [2:0] y_node_1_io_in_0; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 40:26]
  wire [2:0] y_node_1_io_in_2; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 40:26]
  wire [1:0] y_node_1_io_out_0; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 40:26]
  wire [1:0] y_node_1_io_out_2; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 40:26]
  wire [2:0] y_node_2_io_in_0; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 40:26]
  wire [2:0] y_node_2_io_in_2; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 40:26]
  wire [1:0] y_node_2_io_out_0; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 40:26]
  wire [1:0] y_node_2_io_out_2; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 40:26]
  wire [2:0] y_node_3_io_in_0; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 40:26]
  wire [2:0] y_node_3_io_in_2; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 40:26]
  wire [1:0] y_node_3_io_out_0; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 40:26]
  wire [1:0] y_node_3_io_out_2; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 40:26]
  wire [2:0] y_node_4_io_in_0; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 40:26]
  wire [2:0] y_node_4_io_in_2; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 40:26]
  wire [1:0] y_node_4_io_out_0; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 40:26]
  wire [1:0] y_node_4_io_out_2; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 40:26]
  wire [2:0] y_node_5_io_in_0; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 40:26]
  wire [2:0] y_node_5_io_in_2; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 40:26]
  wire [1:0] y_node_5_io_out_0; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 40:26]
  wire [1:0] y_node_5_io_out_2; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 40:26]
  wire [2:0] y_node_6_io_in_0; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 40:26]
  wire [2:0] y_node_6_io_in_2; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 40:26]
  wire [1:0] y_node_6_io_out_0; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 40:26]
  wire [1:0] y_node_6_io_out_2; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 40:26]
  wire [2:0] y_node0_1_io_in_0; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 31:23]
  wire [2:0] y_node0_1_io_in_2; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 31:23]
  wire [1:0] y_node0_1_io_out_0; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 31:23]
  wire [1:0] y_node0_1_io_out_2; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 31:23]
  wire [2:0] y_node_7_io_in_0; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 40:26]
  wire [2:0] y_node_7_io_in_2; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 40:26]
  wire [1:0] y_node_7_io_out_0; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 40:26]
  wire [1:0] y_node_7_io_out_2; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 40:26]
  wire [2:0] y_node_8_io_in_0; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 40:26]
  wire [2:0] y_node_8_io_in_2; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 40:26]
  wire [1:0] y_node_8_io_out_0; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 40:26]
  wire [1:0] y_node_8_io_out_2; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 40:26]
  wire [2:0] y_node_9_io_in_0; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 40:26]
  wire [2:0] y_node_9_io_in_2; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 40:26]
  wire [1:0] y_node_9_io_out_0; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 40:26]
  wire [1:0] y_node_9_io_out_2; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 40:26]
  wire [2:0] y_node_10_io_in_0; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 40:26]
  wire [2:0] y_node_10_io_in_2; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 40:26]
  wire [1:0] y_node_10_io_out_0; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 40:26]
  wire [1:0] y_node_10_io_out_2; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 40:26]
  wire [2:0] y_node0_2_io_in_0; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 31:23]
  wire [2:0] y_node0_2_io_in_2; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 31:23]
  wire [1:0] y_node0_2_io_out_0; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 31:23]
  wire [1:0] y_node0_2_io_out_2; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 31:23]
  wire [2:0] y_node_11_io_in_0; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 40:26]
  wire [2:0] y_node_11_io_in_2; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 40:26]
  wire [1:0] y_node_11_io_out_0; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 40:26]
  wire [1:0] y_node_11_io_out_2; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 40:26]
  wire [2:0] y_node_12_io_in_0; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 40:26]
  wire [2:0] y_node_12_io_in_2; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 40:26]
  wire [1:0] y_node_12_io_out_0; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 40:26]
  wire [1:0] y_node_12_io_out_2; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 40:26]
  wire [2:0] y_node_13_io_in_0; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 40:26]
  wire [2:0] y_node_13_io_in_2; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 40:26]
  wire [1:0] y_node_13_io_out_0; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 40:26]
  wire [1:0] y_node_13_io_out_2; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 40:26]
  wire [2:0] y_node0_3_io_in_0; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 31:23]
  wire [2:0] y_node0_3_io_in_2; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 31:23]
  wire [1:0] y_node0_3_io_out_0; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 31:23]
  wire [1:0] y_node0_3_io_out_2; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 31:23]
  wire [2:0] y_node_14_io_in_0; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 40:26]
  wire [2:0] y_node_14_io_in_2; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 40:26]
  wire [1:0] y_node_14_io_out_0; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 40:26]
  wire [1:0] y_node_14_io_out_2; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 40:26]
  wire [2:0] y_node0_4_io_in_0; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 31:23]
  wire [2:0] y_node0_4_io_in_2; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 31:23]
  wire [1:0] y_node0_4_io_out_0; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 31:23]
  wire [1:0] y_node0_4_io_out_2; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 31:23]
  wire [2:0] y_node_15_io_in_0; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 40:26]
  wire [2:0] y_node_15_io_in_2; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 40:26]
  wire [1:0] y_node_15_io_out_0; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 40:26]
  wire [1:0] y_node_15_io_out_2; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 40:26]
  wire [2:0] y_node0_5_io_in_0; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 31:23]
  wire [2:0] y_node0_5_io_in_2; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 31:23]
  wire [1:0] y_node0_5_io_out_0; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 31:23]
  wire [1:0] y_node0_5_io_out_2; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 31:23]
  wire [2:0] y_node0_6_io_in_0; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 31:23]
  wire [2:0] y_node0_6_io_in_2; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 31:23]
  wire [1:0] y_node0_6_io_out_0; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 31:23]
  wire [1:0] y_node0_6_io_out_2; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 31:23]
  wire  _p_0_T_6 = ~io_e[2]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 23:47]
  wire  p_0 = (io_e[1] | io_e[2] & io_g[1] | ~io_e[2] & io_s[1]) & io_g[0]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 23:67]
  wire  n_0 = (io_e[1] | io_e[2] & io_s[1] | _p_0_T_6 & io_g[1]) & io_s[0]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 24:67]
  wire  z_0 = ~(p_0 | n_0); // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 26:13]
  wire  _p_1_T_6 = ~io_e[3]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 23:47]
  wire  p_1 = (io_e[2] | io_e[3] & io_g[2] | ~io_e[3] & io_s[2]) & io_g[1]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 23:67]
  wire  n_1 = (io_e[2] | io_e[3] & io_s[2] | _p_1_T_6 & io_g[2]) & io_s[1]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 24:67]
  wire  z_1 = ~(p_1 | n_1); // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 26:13]
  wire  _p_2_T_6 = ~io_e[4]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 23:47]
  wire  p_2 = (io_e[3] | io_e[4] & io_g[3] | ~io_e[4] & io_s[3]) & io_g[2]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 23:67]
  wire  n_2 = (io_e[3] | io_e[4] & io_s[3] | _p_2_T_6 & io_g[3]) & io_s[2]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 24:67]
  wire  z_2 = ~(p_2 | n_2); // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 26:13]
  wire  _p_3_T_6 = ~io_e[5]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 23:47]
  wire  p_3 = (io_e[4] | io_e[5] & io_g[4] | ~io_e[5] & io_s[4]) & io_g[3]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 23:67]
  wire  n_3 = (io_e[4] | io_e[5] & io_s[4] | _p_3_T_6 & io_g[4]) & io_s[3]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 24:67]
  wire  z_3 = ~(p_3 | n_3); // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 26:13]
  wire  _p_4_T_6 = ~io_e[6]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 23:47]
  wire  p_4 = (io_e[5] | io_e[6] & io_g[5] | ~io_e[6] & io_s[5]) & io_g[4]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 23:67]
  wire  n_4 = (io_e[5] | io_e[6] & io_s[5] | _p_4_T_6 & io_g[5]) & io_s[4]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 24:67]
  wire  z_4 = ~(p_4 | n_4); // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 26:13]
  wire  _p_5_T_6 = ~io_e[7]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 23:47]
  wire  p_5 = (io_e[6] | io_e[7] & io_g[6] | ~io_e[7] & io_s[6]) & io_g[5]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 23:67]
  wire  n_5 = (io_e[6] | io_e[7] & io_s[6] | _p_5_T_6 & io_g[6]) & io_s[5]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 24:67]
  wire  z_5 = ~(p_5 | n_5); // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 26:13]
  wire  _p_6_T_6 = ~io_e[8]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 23:47]
  wire  p_6 = (io_e[7] | io_e[8] & io_g[7] | ~io_e[8] & io_s[7]) & io_g[6]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 23:67]
  wire  n_6 = (io_e[7] | io_e[8] & io_s[7] | _p_6_T_6 & io_g[7]) & io_s[6]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 24:67]
  wire  z_6 = ~(p_6 | n_6); // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 26:13]
  wire  _p_7_T_6 = ~io_e[9]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 23:47]
  wire  p_7 = (io_e[8] | io_e[9] & io_g[8] | ~io_e[9] & io_s[8]) & io_g[7]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 23:67]
  wire  n_7 = (io_e[8] | io_e[9] & io_s[8] | _p_7_T_6 & io_g[8]) & io_s[7]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 24:67]
  wire  z_7 = ~(p_7 | n_7); // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 26:13]
  wire  _p_8_T_6 = ~io_e[10]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 23:47]
  wire  p_8 = (io_e[9] | io_e[10] & io_g[9] | ~io_e[10] & io_s[9]) & io_g[8]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 23:67]
  wire  n_8 = (io_e[9] | io_e[10] & io_s[9] | _p_8_T_6 & io_g[9]) & io_s[8]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 24:67]
  wire  z_8 = ~(p_8 | n_8); // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 26:13]
  wire  _p_9_T_6 = ~io_e[11]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 23:47]
  wire  p_9 = (io_e[10] | io_e[11] & io_g[10] | ~io_e[11] & io_s[10]) & io_g[9]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 23:67]
  wire  n_9 = (io_e[10] | io_e[11] & io_s[10] | _p_9_T_6 & io_g[10]) & io_s[9]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 24:67]
  wire  z_9 = ~(p_9 | n_9); // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 26:13]
  wire  _p_10_T_6 = ~io_e[12]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 23:47]
  wire  p_10 = (io_e[11] | io_e[12] & io_g[11] | ~io_e[12] & io_s[11]) & io_g[10]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 23:67]
  wire  n_10 = (io_e[11] | io_e[12] & io_s[11] | _p_10_T_6 & io_g[11]) & io_s[10]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 24:67]
  wire  z_10 = ~(p_10 | n_10); // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 26:13]
  wire  _p_11_T_6 = ~io_e[13]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 23:47]
  wire  p_11 = (io_e[12] | io_e[13] & io_g[12] | ~io_e[13] & io_s[12]) & io_g[11]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 23:67]
  wire  n_11 = (io_e[12] | io_e[13] & io_s[12] | _p_11_T_6 & io_g[12]) & io_s[11]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 24:67]
  wire  z_11 = ~(p_11 | n_11); // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 26:13]
  wire  _p_12_T_6 = ~io_e[14]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 23:47]
  wire  p_12 = (io_e[13] | io_e[14] & io_g[13] | ~io_e[14] & io_s[13]) & io_g[12]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 23:67]
  wire  n_12 = (io_e[13] | io_e[14] & io_s[13] | _p_12_T_6 & io_g[13]) & io_s[12]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 24:67]
  wire  z_12 = ~(p_12 | n_12); // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 26:13]
  wire  _p_13_T_6 = ~io_e[15]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 23:47]
  wire  p_13 = (io_e[14] | io_e[15] & io_g[14] | ~io_e[15] & io_s[14]) & io_g[13]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 23:67]
  wire  n_13 = (io_e[14] | io_e[15] & io_s[14] | _p_13_T_6 & io_g[14]) & io_s[13]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 24:67]
  wire  z_13 = ~(p_13 | n_13); // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 26:13]
  wire  _p_14_T_6 = ~io_e[16]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 23:47]
  wire  p_14 = (io_e[15] | io_e[16] & io_g[15] | ~io_e[16] & io_s[15]) & io_g[14]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 23:67]
  wire  n_14 = (io_e[15] | io_e[16] & io_s[15] | _p_14_T_6 & io_g[15]) & io_s[14]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 24:67]
  wire  z_14 = ~(p_14 | n_14); // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 26:13]
  wire  _p_15_T_6 = ~io_e[17]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 23:47]
  wire  p_15 = (io_e[16] | io_e[17] & io_g[16] | ~io_e[17] & io_s[16]) & io_g[15]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 23:67]
  wire  n_15 = (io_e[16] | io_e[17] & io_s[16] | _p_15_T_6 & io_g[16]) & io_s[15]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 24:67]
  wire  z_15 = ~(p_15 | n_15); // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 26:13]
  wire  _p_16_T_6 = ~io_e[18]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 23:47]
  wire  p_16 = (io_e[17] | io_e[18] & io_g[17] | ~io_e[18] & io_s[17]) & io_g[16]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 23:67]
  wire  n_16 = (io_e[17] | io_e[18] & io_s[17] | _p_16_T_6 & io_g[17]) & io_s[16]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 24:67]
  wire  z_16 = ~(p_16 | n_16); // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 26:13]
  wire  _p_17_T_6 = ~io_e[19]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 23:47]
  wire  p_17 = (io_e[18] | io_e[19] & io_g[18] | ~io_e[19] & io_s[18]) & io_g[17]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 23:67]
  wire  n_17 = (io_e[18] | io_e[19] & io_s[18] | _p_17_T_6 & io_g[18]) & io_s[17]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 24:67]
  wire  z_17 = ~(p_17 | n_17); // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 26:13]
  wire  _p_18_T_6 = ~io_e[20]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 23:47]
  wire  p_18 = (io_e[19] | io_e[20] & io_g[19] | ~io_e[20] & io_s[19]) & io_g[18]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 23:67]
  wire  n_18 = (io_e[19] | io_e[20] & io_s[19] | _p_18_T_6 & io_g[19]) & io_s[18]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 24:67]
  wire  z_18 = ~(p_18 | n_18); // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 26:13]
  wire  _p_19_T_6 = ~io_e[21]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 23:47]
  wire  p_19 = (io_e[20] | io_e[21] & io_g[20] | ~io_e[21] & io_s[20]) & io_g[19]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 23:67]
  wire  n_19 = (io_e[20] | io_e[21] & io_s[20] | _p_19_T_6 & io_g[20]) & io_s[19]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 24:67]
  wire  z_19 = ~(p_19 | n_19); // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 26:13]
  wire  _p_20_T_6 = ~io_e[22]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 23:47]
  wire  p_20 = (io_e[21] | io_e[22] & io_g[21] | ~io_e[22] & io_s[21]) & io_g[20]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 23:67]
  wire  n_20 = (io_e[21] | io_e[22] & io_s[21] | _p_20_T_6 & io_g[21]) & io_s[20]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 24:67]
  wire  z_20 = ~(p_20 | n_20); // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 26:13]
  wire  _p_21_T_6 = ~io_e[23]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 23:47]
  wire  p_21 = (io_e[22] | io_e[23] & io_g[22] | ~io_e[23] & io_s[22]) & io_g[21]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 23:67]
  wire  n_21 = (io_e[22] | io_e[23] & io_s[22] | _p_21_T_6 & io_g[22]) & io_s[21]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 24:67]
  wire  z_21 = ~(p_21 | n_21); // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 26:13]
  wire  _p_22_T_6 = ~io_e[24]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 23:47]
  wire  p_22 = (io_e[23] | io_e[24] & io_g[23] | ~io_e[24] & io_s[23]) & io_g[22]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 23:67]
  wire  n_22 = (io_e[23] | io_e[24] & io_s[23] | _p_22_T_6 & io_g[23]) & io_s[22]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 24:67]
  wire  z_22 = ~(p_22 | n_22); // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 26:13]
  wire  p_23 = (io_e[24] | io_g[24]) & io_g[23]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 20:33]
  wire  n_23 = (io_e[24] | io_s[24]) & io_s[23]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 21:33]
  wire  z_23 = ~(p_23 | n_23); // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 26:13]
  wire  z_24 = ~(io_g[24] | io_s[24]); // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 26:13]
  wire [5:0] y_lo_lo = {p_19,p_20,p_21,p_22,p_23,io_g[24]}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 63:28]
  wire [11:0] y_lo = {p_13,p_14,p_15,p_16,p_17,p_18,y_lo_lo}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 63:28]
  wire [5:0] y_hi_lo = {p_7,p_8,p_9,p_10,p_11,p_12}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 63:28]
  wire [24:0] _y_T = {p_0,p_1,p_2,p_3,p_4,p_5,p_6,y_hi_lo,y_lo}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 63:28]
  wire [5:0] y_lo_lo_2 = {z_19,z_20,z_21,z_22,z_23,z_24}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 63:44]
  wire [11:0] y_lo_2 = {z_13,z_14,z_15,z_16,z_17,z_18,y_lo_lo_2}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 63:44]
  wire [5:0] y_hi_lo_2 = {z_7,z_8,z_9,z_10,z_11,z_12}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 63:44]
  wire [24:0] _y_T_2 = {z_0,z_1,z_2,z_3,z_4,z_5,z_6,y_hi_lo_2,y_lo_2}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 63:44]
  wire [1:0] y_node0_io_in_0_hi = {_y_T[2],_y_T[1]}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 32:26]
  wire [1:0] y_node0_io_in_2_hi = {_y_T_2[2],_y_T_2[1]}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 34:26]
  wire  y_nextColumn_p_0 = y_node0_io_out_0[0]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 35:40]
  wire  y_nextColumn_p_1 = y_node0_io_out_0[1]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 35:40]
  wire  y_nextColumn_z_0 = y_node0_io_out_2[0]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 37:40]
  wire  y_nextColumn_z_1 = y_node0_io_out_2[1]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 37:40]
  wire [1:0] y_node_io_in_0_hi = {_y_T[5],_y_T[4]}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 41:29]
  wire [1:0] y_node_io_in_2_hi = {_y_T_2[5],_y_T_2[4]}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 43:29]
  wire  y_pout_0 = y_node_io_out_0[0]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 44:35]
  wire  y_pout_1 = y_node_io_out_0[1]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 44:35]
  wire  y_zout_0 = y_node_io_out_2[0]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 46:35]
  wire  y_zout_1 = y_node_io_out_2[1]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 46:35]
  wire [1:0] y_node_io_in_0_hi_1 = {_y_T[8],_y_T[7]}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 41:29]
  wire [1:0] y_node_io_in_2_hi_1 = {_y_T_2[8],_y_T_2[7]}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 43:29]
  wire  y_pout_0_1 = y_node_1_io_out_0[0]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 44:35]
  wire  y_pout_1_1 = y_node_1_io_out_0[1]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 44:35]
  wire  y_zout_0_1 = y_node_1_io_out_2[0]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 46:35]
  wire  y_zout_1_1 = y_node_1_io_out_2[1]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 46:35]
  wire [1:0] y_node_io_in_0_hi_2 = {_y_T[11],_y_T[10]}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 41:29]
  wire [1:0] y_node_io_in_2_hi_2 = {_y_T_2[11],_y_T_2[10]}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 43:29]
  wire  y_pout_0_2 = y_node_2_io_out_0[0]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 44:35]
  wire  y_pout_1_2 = y_node_2_io_out_0[1]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 44:35]
  wire  y_zout_0_2 = y_node_2_io_out_2[0]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 46:35]
  wire  y_zout_1_2 = y_node_2_io_out_2[1]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 46:35]
  wire [1:0] y_node_io_in_0_hi_3 = {_y_T[14],_y_T[13]}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 41:29]
  wire [1:0] y_node_io_in_2_hi_3 = {_y_T_2[14],_y_T_2[13]}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 43:29]
  wire  y_pout_0_3 = y_node_3_io_out_0[0]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 44:35]
  wire  y_pout_1_3 = y_node_3_io_out_0[1]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 44:35]
  wire  y_zout_0_3 = y_node_3_io_out_2[0]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 46:35]
  wire  y_zout_1_3 = y_node_3_io_out_2[1]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 46:35]
  wire [1:0] y_node_io_in_0_hi_4 = {_y_T[17],_y_T[16]}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 41:29]
  wire [1:0] y_node_io_in_2_hi_4 = {_y_T_2[17],_y_T_2[16]}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 43:29]
  wire  y_pout_0_4 = y_node_4_io_out_0[0]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 44:35]
  wire  y_pout_1_4 = y_node_4_io_out_0[1]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 44:35]
  wire  y_zout_0_4 = y_node_4_io_out_2[0]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 46:35]
  wire  y_zout_1_4 = y_node_4_io_out_2[1]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 46:35]
  wire [1:0] y_node_io_in_0_hi_5 = {_y_T[20],_y_T[19]}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 41:29]
  wire [1:0] y_node_io_in_2_hi_5 = {_y_T_2[20],_y_T_2[19]}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 43:29]
  wire  y_pout_0_5 = y_node_5_io_out_0[0]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 44:35]
  wire  y_pout_1_5 = y_node_5_io_out_0[1]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 44:35]
  wire  y_zout_0_5 = y_node_5_io_out_2[0]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 46:35]
  wire  y_zout_1_5 = y_node_5_io_out_2[1]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 46:35]
  wire [1:0] y_node_io_in_0_hi_6 = {_y_T[23],_y_T[22]}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 41:29]
  wire [1:0] y_node_io_in_2_hi_6 = {_y_T_2[23],_y_T_2[22]}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 43:29]
  wire  y_pout_0_6 = y_node_6_io_out_0[0]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 44:35]
  wire  y_pout_1_6 = y_node_6_io_out_0[1]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 44:35]
  wire  y_zout_0_6 = y_node_6_io_out_2[0]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 46:35]
  wire  y_zout_1_6 = y_node_6_io_out_2[1]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 46:35]
  wire [7:0] y_lo_3 = {y_pout_1_2,y_pout_0_2,y_pout_1_1,y_pout_0_1,y_pout_1,y_pout_0,y_nextColumn_p_1,y_nextColumn_p_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 61:33]
  wire [16:0] _y_T_9 = {_y_T[24],y_pout_1_6,y_pout_0_6,y_pout_1_5,y_pout_0_5,y_pout_1_4,y_pout_0_4,y_pout_1_3,y_pout_0_3
    ,y_lo_3}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 61:33]
  wire [7:0] y_lo_5 = {y_zout_1_2,y_zout_0_2,y_zout_1_1,y_zout_0_1,y_zout_1,y_zout_0,y_nextColumn_z_1,y_nextColumn_z_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 61:87]
  wire [16:0] _y_T_11 = {_y_T_2[24],y_zout_1_6,y_zout_0_6,y_zout_1_5,y_zout_0_5,y_zout_1_4,y_zout_0_4,y_zout_1_3,
    y_zout_0_3,y_lo_5}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 61:87]
  wire [1:0] y_node0_io_in_0_hi_1 = {_y_T_9[2],_y_T_9[1]}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 32:26]
  wire [1:0] y_node0_io_in_2_hi_1 = {_y_T_11[2],_y_T_11[1]}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 34:26]
  wire  y_nextColumn_p_0_1 = y_node0_1_io_out_0[0]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 35:40]
  wire  y_nextColumn_p_1_1 = y_node0_1_io_out_0[1]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 35:40]
  wire  y_nextColumn_z_0_1 = y_node0_1_io_out_2[0]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 37:40]
  wire  y_nextColumn_z_1_1 = y_node0_1_io_out_2[1]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 37:40]
  wire [1:0] y_node_io_in_0_hi_7 = {_y_T_9[5],_y_T_9[4]}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 41:29]
  wire [1:0] y_node_io_in_2_hi_7 = {_y_T_11[5],_y_T_11[4]}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 43:29]
  wire  y_pout_0_7 = y_node_7_io_out_0[0]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 44:35]
  wire  y_pout_1_7 = y_node_7_io_out_0[1]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 44:35]
  wire  y_zout_0_7 = y_node_7_io_out_2[0]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 46:35]
  wire  y_zout_1_7 = y_node_7_io_out_2[1]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 46:35]
  wire [1:0] y_node_io_in_0_hi_8 = {_y_T_9[8],_y_T_9[7]}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 41:29]
  wire [1:0] y_node_io_in_2_hi_8 = {_y_T_11[8],_y_T_11[7]}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 43:29]
  wire  y_pout_0_8 = y_node_8_io_out_0[0]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 44:35]
  wire  y_pout_1_8 = y_node_8_io_out_0[1]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 44:35]
  wire  y_zout_0_8 = y_node_8_io_out_2[0]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 46:35]
  wire  y_zout_1_8 = y_node_8_io_out_2[1]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 46:35]
  wire [1:0] y_node_io_in_0_hi_9 = {_y_T_9[11],_y_T_9[10]}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 41:29]
  wire [1:0] y_node_io_in_2_hi_9 = {_y_T_11[11],_y_T_11[10]}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 43:29]
  wire  y_pout_0_9 = y_node_9_io_out_0[0]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 44:35]
  wire  y_pout_1_9 = y_node_9_io_out_0[1]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 44:35]
  wire  y_zout_0_9 = y_node_9_io_out_2[0]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 46:35]
  wire  y_zout_1_9 = y_node_9_io_out_2[1]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 46:35]
  wire [1:0] y_node_io_in_0_hi_10 = {_y_T_9[14],_y_T_9[13]}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 41:29]
  wire [1:0] y_node_io_in_2_hi_10 = {_y_T_11[14],_y_T_11[13]}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 43:29]
  wire  y_pout_0_10 = y_node_10_io_out_0[0]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 44:35]
  wire  y_pout_1_10 = y_node_10_io_out_0[1]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 44:35]
  wire  y_zout_0_10 = y_node_10_io_out_2[0]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 46:35]
  wire  y_zout_1_10 = y_node_10_io_out_2[1]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 46:35]
  wire [5:0] y_lo_6 = {y_pout_1_8,y_pout_0_8,y_pout_1_7,y_pout_0_7,y_nextColumn_p_1_1,y_nextColumn_p_0_1}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 61:33]
  wire [11:0] _y_T_24 = {_y_T_9[16],_y_T_9[15],y_pout_1_10,y_pout_0_10,y_pout_1_9,y_pout_0_9,y_lo_6}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 61:33]
  wire [5:0] y_lo_8 = {y_zout_1_8,y_zout_0_8,y_zout_1_7,y_zout_0_7,y_nextColumn_z_1_1,y_nextColumn_z_0_1}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 61:87]
  wire [11:0] _y_T_26 = {_y_T_11[16],_y_T_11[15],y_zout_1_10,y_zout_0_10,y_zout_1_9,y_zout_0_9,y_lo_8}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 61:87]
  wire [1:0] y_node0_io_in_0_hi_2 = {_y_T_24[2],_y_T_24[1]}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 32:26]
  wire [1:0] y_node0_io_in_2_hi_2 = {_y_T_26[2],_y_T_26[1]}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 34:26]
  wire  y_nextColumn_p_0_2 = y_node0_2_io_out_0[0]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 35:40]
  wire  y_nextColumn_p_1_2 = y_node0_2_io_out_0[1]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 35:40]
  wire  y_nextColumn_z_0_2 = y_node0_2_io_out_2[0]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 37:40]
  wire  y_nextColumn_z_1_2 = y_node0_2_io_out_2[1]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 37:40]
  wire [1:0] y_node_io_in_0_hi_11 = {_y_T_24[5],_y_T_24[4]}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 41:29]
  wire [1:0] y_node_io_in_2_hi_11 = {_y_T_26[5],_y_T_26[4]}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 43:29]
  wire  y_pout_0_11 = y_node_11_io_out_0[0]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 44:35]
  wire  y_pout_1_11 = y_node_11_io_out_0[1]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 44:35]
  wire  y_zout_0_11 = y_node_11_io_out_2[0]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 46:35]
  wire  y_zout_1_11 = y_node_11_io_out_2[1]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 46:35]
  wire [1:0] y_node_io_in_0_hi_12 = {_y_T_24[8],_y_T_24[7]}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 41:29]
  wire [1:0] y_node_io_in_2_hi_12 = {_y_T_26[8],_y_T_26[7]}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 43:29]
  wire  y_pout_0_12 = y_node_12_io_out_0[0]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 44:35]
  wire  y_pout_1_12 = y_node_12_io_out_0[1]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 44:35]
  wire  y_zout_0_12 = y_node_12_io_out_2[0]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 46:35]
  wire  y_zout_1_12 = y_node_12_io_out_2[1]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 46:35]
  wire [1:0] y_node_io_in_0_hi_13 = {_y_T_24[11],_y_T_24[10]}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 41:29]
  wire [1:0] y_node_io_in_2_hi_13 = {_y_T_26[11],_y_T_26[10]}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 43:29]
  wire  y_pout_0_13 = y_node_13_io_out_0[0]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 44:35]
  wire  y_pout_1_13 = y_node_13_io_out_0[1]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 44:35]
  wire  y_zout_0_13 = y_node_13_io_out_2[0]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 46:35]
  wire  y_zout_1_13 = y_node_13_io_out_2[1]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 46:35]
  wire [7:0] _y_T_27 = {y_pout_1_13,y_pout_0_13,y_pout_1_12,y_pout_0_12,y_pout_1_11,y_pout_0_11,y_nextColumn_p_1_2,
    y_nextColumn_p_0_2}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 61:33]
  wire [7:0] _y_T_29 = {y_zout_1_13,y_zout_0_13,y_zout_1_12,y_zout_0_12,y_zout_1_11,y_zout_0_11,y_nextColumn_z_1_2,
    y_nextColumn_z_0_2}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 61:87]
  wire [1:0] y_node0_io_in_0_hi_3 = {_y_T_27[2],_y_T_27[1]}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 32:26]
  wire [1:0] y_node0_io_in_2_hi_3 = {_y_T_29[2],_y_T_29[1]}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 34:26]
  wire  y_nextColumn_p_0_3 = y_node0_3_io_out_0[0]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 35:40]
  wire  y_nextColumn_p_1_3 = y_node0_3_io_out_0[1]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 35:40]
  wire  y_nextColumn_z_0_3 = y_node0_3_io_out_2[0]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 37:40]
  wire  y_nextColumn_z_1_3 = y_node0_3_io_out_2[1]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 37:40]
  wire [1:0] y_node_io_in_0_hi_14 = {_y_T_27[5],_y_T_27[4]}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 41:29]
  wire [1:0] y_node_io_in_2_hi_14 = {_y_T_29[5],_y_T_29[4]}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 43:29]
  wire  y_pout_0_14 = y_node_14_io_out_0[0]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 44:35]
  wire  y_pout_1_14 = y_node_14_io_out_0[1]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 44:35]
  wire  y_zout_0_14 = y_node_14_io_out_2[0]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 46:35]
  wire  y_zout_1_14 = y_node_14_io_out_2[1]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 46:35]
  wire [5:0] _y_T_42 = {_y_T_27[7],_y_T_27[6],y_pout_1_14,y_pout_0_14,y_nextColumn_p_1_3,y_nextColumn_p_0_3}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 61:33]
  wire [5:0] _y_T_44 = {_y_T_29[7],_y_T_29[6],y_zout_1_14,y_zout_0_14,y_nextColumn_z_1_3,y_nextColumn_z_0_3}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 61:87]
  wire [1:0] y_node0_io_in_0_hi_4 = {_y_T_42[2],_y_T_42[1]}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 32:26]
  wire [1:0] y_node0_io_in_2_hi_4 = {_y_T_44[2],_y_T_44[1]}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 34:26]
  wire  y_nextColumn_p_0_4 = y_node0_4_io_out_0[0]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 35:40]
  wire  y_nextColumn_p_1_4 = y_node0_4_io_out_0[1]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 35:40]
  wire  y_nextColumn_z_0_4 = y_node0_4_io_out_2[0]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 37:40]
  wire  y_nextColumn_z_1_4 = y_node0_4_io_out_2[1]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 37:40]
  wire [1:0] y_node_io_in_0_hi_15 = {_y_T_42[5],_y_T_42[4]}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 41:29]
  wire [1:0] y_node_io_in_2_hi_15 = {_y_T_44[5],_y_T_44[4]}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 43:29]
  wire  y_pout_0_15 = y_node_15_io_out_0[0]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 44:35]
  wire  y_pout_1_15 = y_node_15_io_out_0[1]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 44:35]
  wire  y_zout_0_15 = y_node_15_io_out_2[0]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 46:35]
  wire  y_zout_1_15 = y_node_15_io_out_2[1]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 46:35]
  wire [3:0] _y_T_45 = {y_pout_1_15,y_pout_0_15,y_nextColumn_p_1_4,y_nextColumn_p_0_4}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 61:33]
  wire [3:0] _y_T_47 = {y_zout_1_15,y_zout_0_15,y_nextColumn_z_1_4,y_nextColumn_z_0_4}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 61:87]
  wire [1:0] y_node0_io_in_0_hi_5 = {_y_T_45[2],_y_T_45[1]}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 32:26]
  wire [1:0] y_node0_io_in_2_hi_5 = {_y_T_47[2],_y_T_47[1]}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 34:26]
  wire  y_nextColumn_p_0_5 = y_node0_5_io_out_0[0]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 35:40]
  wire  y_nextColumn_p_1_5 = y_node0_5_io_out_0[1]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 35:40]
  wire  y_nextColumn_z_0_5 = y_node0_5_io_out_2[0]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 37:40]
  wire  y_nextColumn_z_1_5 = y_node0_5_io_out_2[1]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 37:40]
  wire [2:0] _y_T_54 = {_y_T_45[3],y_nextColumn_p_1_5,y_nextColumn_p_0_5}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 61:33]
  wire [2:0] _y_T_56 = {_y_T_47[3],y_nextColumn_z_1_5,y_nextColumn_z_0_5}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 61:87]
  wire [1:0] y_node0_io_in_0_hi_6 = {_y_T_54[2],_y_T_54[1]}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 32:26]
  wire [1:0] y_node0_io_in_2_hi_6 = {_y_T_56[2],_y_T_56[1]}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 34:26]
  wire  y_nextColumn_p_0_6 = y_node0_6_io_out_0[0]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 35:40]
  wire  y_nextColumn_p_1_6 = y_node0_6_io_out_0[1]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 35:40]
  wire  y_nextColumn_z_0_6 = y_node0_6_io_out_2[0]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 37:40]
  wire  y_nextColumn_z_1_6 = y_node0_6_io_out_2[1]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 37:40]
  node y_node0 ( // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 31:23]
    .io_in_0(y_node0_io_in_0),
    .io_in_2(y_node0_io_in_2),
    .io_out_0(y_node0_io_out_0),
    .io_out_2(y_node0_io_out_2)
  );
  node y_node ( // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 40:26]
    .io_in_0(y_node_io_in_0),
    .io_in_2(y_node_io_in_2),
    .io_out_0(y_node_io_out_0),
    .io_out_2(y_node_io_out_2)
  );
  node y_node_1 ( // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 40:26]
    .io_in_0(y_node_1_io_in_0),
    .io_in_2(y_node_1_io_in_2),
    .io_out_0(y_node_1_io_out_0),
    .io_out_2(y_node_1_io_out_2)
  );
  node y_node_2 ( // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 40:26]
    .io_in_0(y_node_2_io_in_0),
    .io_in_2(y_node_2_io_in_2),
    .io_out_0(y_node_2_io_out_0),
    .io_out_2(y_node_2_io_out_2)
  );
  node y_node_3 ( // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 40:26]
    .io_in_0(y_node_3_io_in_0),
    .io_in_2(y_node_3_io_in_2),
    .io_out_0(y_node_3_io_out_0),
    .io_out_2(y_node_3_io_out_2)
  );
  node y_node_4 ( // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 40:26]
    .io_in_0(y_node_4_io_in_0),
    .io_in_2(y_node_4_io_in_2),
    .io_out_0(y_node_4_io_out_0),
    .io_out_2(y_node_4_io_out_2)
  );
  node y_node_5 ( // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 40:26]
    .io_in_0(y_node_5_io_in_0),
    .io_in_2(y_node_5_io_in_2),
    .io_out_0(y_node_5_io_out_0),
    .io_out_2(y_node_5_io_out_2)
  );
  node y_node_6 ( // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 40:26]
    .io_in_0(y_node_6_io_in_0),
    .io_in_2(y_node_6_io_in_2),
    .io_out_0(y_node_6_io_out_0),
    .io_out_2(y_node_6_io_out_2)
  );
  node y_node0_1 ( // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 31:23]
    .io_in_0(y_node0_1_io_in_0),
    .io_in_2(y_node0_1_io_in_2),
    .io_out_0(y_node0_1_io_out_0),
    .io_out_2(y_node0_1_io_out_2)
  );
  node y_node_7 ( // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 40:26]
    .io_in_0(y_node_7_io_in_0),
    .io_in_2(y_node_7_io_in_2),
    .io_out_0(y_node_7_io_out_0),
    .io_out_2(y_node_7_io_out_2)
  );
  node y_node_8 ( // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 40:26]
    .io_in_0(y_node_8_io_in_0),
    .io_in_2(y_node_8_io_in_2),
    .io_out_0(y_node_8_io_out_0),
    .io_out_2(y_node_8_io_out_2)
  );
  node y_node_9 ( // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 40:26]
    .io_in_0(y_node_9_io_in_0),
    .io_in_2(y_node_9_io_in_2),
    .io_out_0(y_node_9_io_out_0),
    .io_out_2(y_node_9_io_out_2)
  );
  node y_node_10 ( // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 40:26]
    .io_in_0(y_node_10_io_in_0),
    .io_in_2(y_node_10_io_in_2),
    .io_out_0(y_node_10_io_out_0),
    .io_out_2(y_node_10_io_out_2)
  );
  node y_node0_2 ( // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 31:23]
    .io_in_0(y_node0_2_io_in_0),
    .io_in_2(y_node0_2_io_in_2),
    .io_out_0(y_node0_2_io_out_0),
    .io_out_2(y_node0_2_io_out_2)
  );
  node y_node_11 ( // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 40:26]
    .io_in_0(y_node_11_io_in_0),
    .io_in_2(y_node_11_io_in_2),
    .io_out_0(y_node_11_io_out_0),
    .io_out_2(y_node_11_io_out_2)
  );
  node y_node_12 ( // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 40:26]
    .io_in_0(y_node_12_io_in_0),
    .io_in_2(y_node_12_io_in_2),
    .io_out_0(y_node_12_io_out_0),
    .io_out_2(y_node_12_io_out_2)
  );
  node y_node_13 ( // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 40:26]
    .io_in_0(y_node_13_io_in_0),
    .io_in_2(y_node_13_io_in_2),
    .io_out_0(y_node_13_io_out_0),
    .io_out_2(y_node_13_io_out_2)
  );
  node y_node0_3 ( // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 31:23]
    .io_in_0(y_node0_3_io_in_0),
    .io_in_2(y_node0_3_io_in_2),
    .io_out_0(y_node0_3_io_out_0),
    .io_out_2(y_node0_3_io_out_2)
  );
  node y_node_14 ( // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 40:26]
    .io_in_0(y_node_14_io_in_0),
    .io_in_2(y_node_14_io_in_2),
    .io_out_0(y_node_14_io_out_0),
    .io_out_2(y_node_14_io_out_2)
  );
  node y_node0_4 ( // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 31:23]
    .io_in_0(y_node0_4_io_in_0),
    .io_in_2(y_node0_4_io_in_2),
    .io_out_0(y_node0_4_io_out_0),
    .io_out_2(y_node0_4_io_out_2)
  );
  node y_node_15 ( // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 40:26]
    .io_in_0(y_node_15_io_in_0),
    .io_in_2(y_node_15_io_in_2),
    .io_out_0(y_node_15_io_out_0),
    .io_out_2(y_node_15_io_out_2)
  );
  node y_node0_5 ( // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 31:23]
    .io_in_0(y_node0_5_io_in_0),
    .io_in_2(y_node0_5_io_in_2),
    .io_out_0(y_node0_5_io_out_0),
    .io_out_2(y_node0_5_io_out_2)
  );
  node y_node0_6 ( // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 31:23]
    .io_in_0(y_node0_6_io_in_0),
    .io_in_2(y_node0_6_io_in_2),
    .io_out_0(y_node0_6_io_out_0),
    .io_out_2(y_node0_6_io_out_2)
  );
  assign io_y = (y_nextColumn_p_0_6 ^ y_nextColumn_p_1_6) & ~y_nextColumn_z_0_6 & ~y_nextColumn_z_1_6; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 60:81]
  assign y_node0_io_in_0 = {y_node0_io_in_0_hi,_y_T[0]}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 32:26]
  assign y_node0_io_in_2 = {y_node0_io_in_2_hi,_y_T_2[0]}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 34:26]
  assign y_node_io_in_0 = {y_node_io_in_0_hi,_y_T[3]}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 41:29]
  assign y_node_io_in_2 = {y_node_io_in_2_hi,_y_T_2[3]}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 43:29]
  assign y_node_1_io_in_0 = {y_node_io_in_0_hi_1,_y_T[6]}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 41:29]
  assign y_node_1_io_in_2 = {y_node_io_in_2_hi_1,_y_T_2[6]}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 43:29]
  assign y_node_2_io_in_0 = {y_node_io_in_0_hi_2,_y_T[9]}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 41:29]
  assign y_node_2_io_in_2 = {y_node_io_in_2_hi_2,_y_T_2[9]}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 43:29]
  assign y_node_3_io_in_0 = {y_node_io_in_0_hi_3,_y_T[12]}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 41:29]
  assign y_node_3_io_in_2 = {y_node_io_in_2_hi_3,_y_T_2[12]}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 43:29]
  assign y_node_4_io_in_0 = {y_node_io_in_0_hi_4,_y_T[15]}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 41:29]
  assign y_node_4_io_in_2 = {y_node_io_in_2_hi_4,_y_T_2[15]}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 43:29]
  assign y_node_5_io_in_0 = {y_node_io_in_0_hi_5,_y_T[18]}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 41:29]
  assign y_node_5_io_in_2 = {y_node_io_in_2_hi_5,_y_T_2[18]}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 43:29]
  assign y_node_6_io_in_0 = {y_node_io_in_0_hi_6,_y_T[21]}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 41:29]
  assign y_node_6_io_in_2 = {y_node_io_in_2_hi_6,_y_T_2[21]}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 43:29]
  assign y_node0_1_io_in_0 = {y_node0_io_in_0_hi_1,_y_T_9[0]}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 32:26]
  assign y_node0_1_io_in_2 = {y_node0_io_in_2_hi_1,_y_T_11[0]}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 34:26]
  assign y_node_7_io_in_0 = {y_node_io_in_0_hi_7,_y_T_9[3]}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 41:29]
  assign y_node_7_io_in_2 = {y_node_io_in_2_hi_7,_y_T_11[3]}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 43:29]
  assign y_node_8_io_in_0 = {y_node_io_in_0_hi_8,_y_T_9[6]}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 41:29]
  assign y_node_8_io_in_2 = {y_node_io_in_2_hi_8,_y_T_11[6]}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 43:29]
  assign y_node_9_io_in_0 = {y_node_io_in_0_hi_9,_y_T_9[9]}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 41:29]
  assign y_node_9_io_in_2 = {y_node_io_in_2_hi_9,_y_T_11[9]}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 43:29]
  assign y_node_10_io_in_0 = {y_node_io_in_0_hi_10,_y_T_9[12]}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 41:29]
  assign y_node_10_io_in_2 = {y_node_io_in_2_hi_10,_y_T_11[12]}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 43:29]
  assign y_node0_2_io_in_0 = {y_node0_io_in_0_hi_2,_y_T_24[0]}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 32:26]
  assign y_node0_2_io_in_2 = {y_node0_io_in_2_hi_2,_y_T_26[0]}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 34:26]
  assign y_node_11_io_in_0 = {y_node_io_in_0_hi_11,_y_T_24[3]}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 41:29]
  assign y_node_11_io_in_2 = {y_node_io_in_2_hi_11,_y_T_26[3]}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 43:29]
  assign y_node_12_io_in_0 = {y_node_io_in_0_hi_12,_y_T_24[6]}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 41:29]
  assign y_node_12_io_in_2 = {y_node_io_in_2_hi_12,_y_T_26[6]}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 43:29]
  assign y_node_13_io_in_0 = {y_node_io_in_0_hi_13,_y_T_24[9]}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 41:29]
  assign y_node_13_io_in_2 = {y_node_io_in_2_hi_13,_y_T_26[9]}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 43:29]
  assign y_node0_3_io_in_0 = {y_node0_io_in_0_hi_3,_y_T_27[0]}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 32:26]
  assign y_node0_3_io_in_2 = {y_node0_io_in_2_hi_3,_y_T_29[0]}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 34:26]
  assign y_node_14_io_in_0 = {y_node_io_in_0_hi_14,_y_T_27[3]}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 41:29]
  assign y_node_14_io_in_2 = {y_node_io_in_2_hi_14,_y_T_29[3]}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 43:29]
  assign y_node0_4_io_in_0 = {y_node0_io_in_0_hi_4,_y_T_42[0]}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 32:26]
  assign y_node0_4_io_in_2 = {y_node0_io_in_2_hi_4,_y_T_44[0]}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 34:26]
  assign y_node_15_io_in_0 = {y_node_io_in_0_hi_15,_y_T_42[3]}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 41:29]
  assign y_node_15_io_in_2 = {y_node_io_in_2_hi_15,_y_T_44[3]}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 43:29]
  assign y_node0_5_io_in_0 = {y_node0_io_in_0_hi_5,_y_T_45[0]}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 32:26]
  assign y_node0_5_io_in_2 = {y_node0_io_in_2_hi_5,_y_T_47[0]}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 34:26]
  assign y_node0_6_io_in_0 = {y_node0_io_in_0_hi_6,_y_T_54[0]}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 32:26]
  assign y_node0_6_io_in_2 = {y_node0_io_in_2_hi_6,_y_T_56[0]}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/ErrorDetector.scala 34:26]
endmodule
module LZC_9(
  input  [24:0] io_in, // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/LZC.scala 11:14]
  output [4:0]  io_out // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/LZC.scala 11:14]
);
  wire [4:0] _io_out_T_25 = io_in[1] ? 5'h17 : 5'h18; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [4:0] _io_out_T_26 = io_in[2] ? 5'h16 : _io_out_T_25; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [4:0] _io_out_T_27 = io_in[3] ? 5'h15 : _io_out_T_26; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [4:0] _io_out_T_28 = io_in[4] ? 5'h14 : _io_out_T_27; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [4:0] _io_out_T_29 = io_in[5] ? 5'h13 : _io_out_T_28; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [4:0] _io_out_T_30 = io_in[6] ? 5'h12 : _io_out_T_29; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [4:0] _io_out_T_31 = io_in[7] ? 5'h11 : _io_out_T_30; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [4:0] _io_out_T_32 = io_in[8] ? 5'h10 : _io_out_T_31; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [4:0] _io_out_T_33 = io_in[9] ? 5'hf : _io_out_T_32; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [4:0] _io_out_T_34 = io_in[10] ? 5'he : _io_out_T_33; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [4:0] _io_out_T_35 = io_in[11] ? 5'hd : _io_out_T_34; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [4:0] _io_out_T_36 = io_in[12] ? 5'hc : _io_out_T_35; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [4:0] _io_out_T_37 = io_in[13] ? 5'hb : _io_out_T_36; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [4:0] _io_out_T_38 = io_in[14] ? 5'ha : _io_out_T_37; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [4:0] _io_out_T_39 = io_in[15] ? 5'h9 : _io_out_T_38; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [4:0] _io_out_T_40 = io_in[16] ? 5'h8 : _io_out_T_39; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [4:0] _io_out_T_41 = io_in[17] ? 5'h7 : _io_out_T_40; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [4:0] _io_out_T_42 = io_in[18] ? 5'h6 : _io_out_T_41; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [4:0] _io_out_T_43 = io_in[19] ? 5'h5 : _io_out_T_42; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [4:0] _io_out_T_44 = io_in[20] ? 5'h4 : _io_out_T_43; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [4:0] _io_out_T_45 = io_in[21] ? 5'h3 : _io_out_T_44; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [4:0] _io_out_T_46 = io_in[22] ? 5'h2 : _io_out_T_45; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [4:0] _io_out_T_47 = io_in[23] ? 5'h1 : _io_out_T_46; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  assign io_out = io_in[24] ? 5'h0 : _io_out_T_47; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
endmodule
module LZA(
  input  [24:0] io_a, // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/LZA.scala 15:14]
  input  [24:0] io_b, // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/LZA.scala 15:14]
  output [4:0]  io_lzc, // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/LZA.scala 15:14]
  output        io_error, // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/LZA.scala 15:14]
  output        io_zero // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/LZA.scala 15:14]
);
  wire [24:0] preEncoder_io_g; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/LZA.scala 24:26]
  wire [24:0] preEncoder_io_s; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/LZA.scala 24:26]
  wire [24:0] preEncoder_io_e; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/LZA.scala 24:26]
  wire [24:0] preEncoder_io_f; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/LZA.scala 24:26]
  wire [24:0] errorDetector_io_g; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/LZA.scala 30:29]
  wire [24:0] errorDetector_io_s; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/LZA.scala 30:29]
  wire [24:0] errorDetector_io_e; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/LZA.scala 30:29]
  wire  errorDetector_io_y; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/LZA.scala 30:29]
  wire [24:0] io_lzc_lzc_io_in; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/LZC.scala 21:21]
  wire [4:0] io_lzc_lzc_io_out; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/LZC.scala 21:21]
  wire  g_0 = io_a[0] & ~io_b[0]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/LZA.scala 19:18]
  wire  s_0 = ~io_a[0] & io_b[0]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/LZA.scala 20:21]
  wire  e_0 = ~(io_a[0] ^ io_b[0]); // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/LZA.scala 21:13]
  wire  g_1 = io_a[1] & ~io_b[1]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/LZA.scala 19:18]
  wire  s_1 = ~io_a[1] & io_b[1]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/LZA.scala 20:21]
  wire  e_1 = ~(io_a[1] ^ io_b[1]); // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/LZA.scala 21:13]
  wire  g_2 = io_a[2] & ~io_b[2]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/LZA.scala 19:18]
  wire  s_2 = ~io_a[2] & io_b[2]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/LZA.scala 20:21]
  wire  e_2 = ~(io_a[2] ^ io_b[2]); // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/LZA.scala 21:13]
  wire  g_3 = io_a[3] & ~io_b[3]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/LZA.scala 19:18]
  wire  s_3 = ~io_a[3] & io_b[3]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/LZA.scala 20:21]
  wire  e_3 = ~(io_a[3] ^ io_b[3]); // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/LZA.scala 21:13]
  wire  g_4 = io_a[4] & ~io_b[4]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/LZA.scala 19:18]
  wire  s_4 = ~io_a[4] & io_b[4]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/LZA.scala 20:21]
  wire  e_4 = ~(io_a[4] ^ io_b[4]); // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/LZA.scala 21:13]
  wire  g_5 = io_a[5] & ~io_b[5]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/LZA.scala 19:18]
  wire  s_5 = ~io_a[5] & io_b[5]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/LZA.scala 20:21]
  wire  e_5 = ~(io_a[5] ^ io_b[5]); // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/LZA.scala 21:13]
  wire  g_6 = io_a[6] & ~io_b[6]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/LZA.scala 19:18]
  wire  s_6 = ~io_a[6] & io_b[6]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/LZA.scala 20:21]
  wire  e_6 = ~(io_a[6] ^ io_b[6]); // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/LZA.scala 21:13]
  wire  g_7 = io_a[7] & ~io_b[7]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/LZA.scala 19:18]
  wire  s_7 = ~io_a[7] & io_b[7]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/LZA.scala 20:21]
  wire  e_7 = ~(io_a[7] ^ io_b[7]); // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/LZA.scala 21:13]
  wire  g_8 = io_a[8] & ~io_b[8]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/LZA.scala 19:18]
  wire  s_8 = ~io_a[8] & io_b[8]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/LZA.scala 20:21]
  wire  e_8 = ~(io_a[8] ^ io_b[8]); // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/LZA.scala 21:13]
  wire  g_9 = io_a[9] & ~io_b[9]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/LZA.scala 19:18]
  wire  s_9 = ~io_a[9] & io_b[9]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/LZA.scala 20:21]
  wire  e_9 = ~(io_a[9] ^ io_b[9]); // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/LZA.scala 21:13]
  wire  g_10 = io_a[10] & ~io_b[10]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/LZA.scala 19:18]
  wire  s_10 = ~io_a[10] & io_b[10]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/LZA.scala 20:21]
  wire  e_10 = ~(io_a[10] ^ io_b[10]); // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/LZA.scala 21:13]
  wire  g_11 = io_a[11] & ~io_b[11]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/LZA.scala 19:18]
  wire  s_11 = ~io_a[11] & io_b[11]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/LZA.scala 20:21]
  wire  e_11 = ~(io_a[11] ^ io_b[11]); // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/LZA.scala 21:13]
  wire  g_12 = io_a[12] & ~io_b[12]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/LZA.scala 19:18]
  wire  s_12 = ~io_a[12] & io_b[12]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/LZA.scala 20:21]
  wire  e_12 = ~(io_a[12] ^ io_b[12]); // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/LZA.scala 21:13]
  wire  g_13 = io_a[13] & ~io_b[13]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/LZA.scala 19:18]
  wire  s_13 = ~io_a[13] & io_b[13]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/LZA.scala 20:21]
  wire  e_13 = ~(io_a[13] ^ io_b[13]); // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/LZA.scala 21:13]
  wire  g_14 = io_a[14] & ~io_b[14]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/LZA.scala 19:18]
  wire  s_14 = ~io_a[14] & io_b[14]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/LZA.scala 20:21]
  wire  e_14 = ~(io_a[14] ^ io_b[14]); // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/LZA.scala 21:13]
  wire  g_15 = io_a[15] & ~io_b[15]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/LZA.scala 19:18]
  wire  s_15 = ~io_a[15] & io_b[15]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/LZA.scala 20:21]
  wire  e_15 = ~(io_a[15] ^ io_b[15]); // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/LZA.scala 21:13]
  wire  g_16 = io_a[16] & ~io_b[16]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/LZA.scala 19:18]
  wire  s_16 = ~io_a[16] & io_b[16]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/LZA.scala 20:21]
  wire  e_16 = ~(io_a[16] ^ io_b[16]); // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/LZA.scala 21:13]
  wire  g_17 = io_a[17] & ~io_b[17]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/LZA.scala 19:18]
  wire  s_17 = ~io_a[17] & io_b[17]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/LZA.scala 20:21]
  wire  e_17 = ~(io_a[17] ^ io_b[17]); // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/LZA.scala 21:13]
  wire  g_18 = io_a[18] & ~io_b[18]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/LZA.scala 19:18]
  wire  s_18 = ~io_a[18] & io_b[18]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/LZA.scala 20:21]
  wire  e_18 = ~(io_a[18] ^ io_b[18]); // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/LZA.scala 21:13]
  wire  g_19 = io_a[19] & ~io_b[19]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/LZA.scala 19:18]
  wire  s_19 = ~io_a[19] & io_b[19]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/LZA.scala 20:21]
  wire  e_19 = ~(io_a[19] ^ io_b[19]); // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/LZA.scala 21:13]
  wire  g_20 = io_a[20] & ~io_b[20]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/LZA.scala 19:18]
  wire  s_20 = ~io_a[20] & io_b[20]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/LZA.scala 20:21]
  wire  e_20 = ~(io_a[20] ^ io_b[20]); // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/LZA.scala 21:13]
  wire  g_21 = io_a[21] & ~io_b[21]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/LZA.scala 19:18]
  wire  s_21 = ~io_a[21] & io_b[21]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/LZA.scala 20:21]
  wire  e_21 = ~(io_a[21] ^ io_b[21]); // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/LZA.scala 21:13]
  wire  g_22 = io_a[22] & ~io_b[22]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/LZA.scala 19:18]
  wire  s_22 = ~io_a[22] & io_b[22]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/LZA.scala 20:21]
  wire  e_22 = ~(io_a[22] ^ io_b[22]); // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/LZA.scala 21:13]
  wire  g_23 = io_a[23] & ~io_b[23]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/LZA.scala 19:18]
  wire  s_23 = ~io_a[23] & io_b[23]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/LZA.scala 20:21]
  wire  e_23 = ~(io_a[23] ^ io_b[23]); // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/LZA.scala 21:13]
  wire  g_24 = io_a[24] & ~io_b[24]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/LZA.scala 19:18]
  wire  s_24 = ~io_a[24] & io_b[24]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/LZA.scala 20:21]
  wire  e_24 = ~(io_a[24] ^ io_b[24]); // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/LZA.scala 21:13]
  wire [5:0] preEncoder_io_g_lo_lo = {g_5,g_4,g_3,g_2,g_1,g_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/LZA.scala 25:25]
  wire [11:0] preEncoder_io_g_lo = {g_11,g_10,g_9,g_8,g_7,g_6,preEncoder_io_g_lo_lo}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/LZA.scala 25:25]
  wire [5:0] preEncoder_io_g_hi_lo = {g_17,g_16,g_15,g_14,g_13,g_12}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/LZA.scala 25:25]
  wire [12:0] preEncoder_io_g_hi = {g_24,g_23,g_22,g_21,g_20,g_19,g_18,preEncoder_io_g_hi_lo}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/LZA.scala 25:25]
  wire [5:0] preEncoder_io_s_lo_lo = {s_5,s_4,s_3,s_2,s_1,s_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/LZA.scala 26:25]
  wire [11:0] preEncoder_io_s_lo = {s_11,s_10,s_9,s_8,s_7,s_6,preEncoder_io_s_lo_lo}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/LZA.scala 26:25]
  wire [5:0] preEncoder_io_s_hi_lo = {s_17,s_16,s_15,s_14,s_13,s_12}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/LZA.scala 26:25]
  wire [12:0] preEncoder_io_s_hi = {s_24,s_23,s_22,s_21,s_20,s_19,s_18,preEncoder_io_s_hi_lo}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/LZA.scala 26:25]
  wire [5:0] preEncoder_io_e_lo_lo = {e_5,e_4,e_3,e_2,e_1,e_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/LZA.scala 27:25]
  wire [11:0] preEncoder_io_e_lo = {e_11,e_10,e_9,e_8,e_7,e_6,preEncoder_io_e_lo_lo}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/LZA.scala 27:25]
  wire [5:0] preEncoder_io_e_hi_lo = {e_17,e_16,e_15,e_14,e_13,e_12}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/LZA.scala 27:25]
  wire [12:0] preEncoder_io_e_hi = {e_24,e_23,e_22,e_21,e_20,e_19,e_18,preEncoder_io_e_hi_lo}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/LZA.scala 27:25]
  PreEncoder preEncoder ( // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/LZA.scala 24:26]
    .io_g(preEncoder_io_g),
    .io_s(preEncoder_io_s),
    .io_e(preEncoder_io_e),
    .io_f(preEncoder_io_f)
  );
  ErrorDetector errorDetector ( // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/LZA.scala 30:29]
    .io_g(errorDetector_io_g),
    .io_s(errorDetector_io_s),
    .io_e(errorDetector_io_e),
    .io_y(errorDetector_io_y)
  );
  LZC_9 io_lzc_lzc ( // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/LZC.scala 21:21]
    .io_in(io_lzc_lzc_io_in),
    .io_out(io_lzc_lzc_io_out)
  );
  assign io_lzc = io_lzc_lzc_io_out; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/LZA.scala 36:10]
  assign io_error = errorDetector_io_y; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/LZA.scala 35:12]
  assign io_zero = ~(|preEncoder_io_f); // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/LZA.scala 37:14]
  assign preEncoder_io_g = {preEncoder_io_g_hi,preEncoder_io_g_lo}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/LZA.scala 25:25]
  assign preEncoder_io_s = {preEncoder_io_s_hi,preEncoder_io_s_lo}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/LZA.scala 26:25]
  assign preEncoder_io_e = {preEncoder_io_e_hi,preEncoder_io_e_lo}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/LZA.scala 27:25]
  assign errorDetector_io_g = {preEncoder_io_g_hi,preEncoder_io_g_lo}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/LZA.scala 31:27]
  assign errorDetector_io_s = {preEncoder_io_s_hi,preEncoder_io_s_lo}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/LZA.scala 32:27]
  assign errorDetector_io_e = {preEncoder_io_e_hi,preEncoder_io_e_lo}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/LZA.scala 33:27]
  assign io_lzc_lzc_io_in = preEncoder_io_f; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/lza_utils/LZC.scala 22:15]
endmodule
module ClosePath(
  input         io_in_a_sign, // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FADD.scala 108:14]
  input  [7:0]  io_in_a_exp, // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FADD.scala 108:14]
  input  [23:0] io_in_a_sig, // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FADD.scala 108:14]
  input  [7:0]  io_in_b_exp, // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FADD.scala 108:14]
  input  [23:0] io_in_b_sig, // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FADD.scala 108:14]
  input         io_in_needShift, // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FADD.scala 108:14]
  output [31:0] io_out_result, // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FADD.scala 108:14]
  output        io_out_near_path_of // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FADD.scala 108:14]
);
  wire [24:0] lza_io_a; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FADD.scala 134:19]
  wire [24:0] lza_io_b; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FADD.scala 134:19]
  wire [4:0] lza_io_lzc; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FADD.scala 134:19]
  wire  lza_io_error; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FADD.scala 134:19]
  wire  lza_io_zero; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FADD.scala 134:19]
  wire [26:0] near_path_tininess_rounder_io_in_sig; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FADD.scala 174:42]
  wire [22:0] near_path_rounder_io_in; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/RoundingUnit.scala 44:25]
  wire  near_path_rounder_io_roundIn; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/RoundingUnit.scala 44:25]
  wire  near_path_rounder_io_stickyIn; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/RoundingUnit.scala 44:25]
  wire [22:0] near_path_rounder_io_out; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/RoundingUnit.scala 44:25]
  wire  near_path_rounder_io_cout; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/RoundingUnit.scala 44:25]
  wire [24:0] _b_sig_T = {io_in_b_sig,1'h0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FADD.scala 123:19]
  wire [24:0] b_sig = _b_sig_T >> io_in_needShift; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FADD.scala 123:43]
  wire  bIsZero = ~(|io_in_b_exp); // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FADD.scala 124:17]
  wire [25:0] _resultSigComplementForm_T = {1'h0,io_in_a_sig,1'h0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FADD.scala 126:8]
  wire [24:0] _resultSigComplementForm_T_2 = ~b_sig; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FADD.scala 127:42]
  wire [24:0] _resultSigComplementForm_T_4 = _resultSigComplementForm_T_2 + 25'h1; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FADD.scala 127:49]
  wire [25:0] _resultSigComplementForm_T_5 = {1'h1,_resultSigComplementForm_T_4}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FADD.scala 127:31]
  wire [25:0] _resultSigComplementForm_T_7 = _resultSigComplementForm_T + _resultSigComplementForm_T_5; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FADD.scala 127:26]
  wire [25:0] resultSigComplementForm = bIsZero ? _resultSigComplementForm_T : _resultSigComplementForm_T_7; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FADD.scala 125:36]
  wire  a_LessThan_b = resultSigComplementForm[25]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FADD.scala 128:50]
  wire [24:0] _resultSigNoRound_T_1 = ~resultSigComplementForm[24:0]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FADD.scala 130:5]
  wire [24:0] _resultSigNoRound_T_3 = _resultSigNoRound_T_1 + 25'h1; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FADD.scala 130:38]
  wire [24:0] resultSigNoRound = a_LessThan_b ? _resultSigNoRound_T_3 : resultSigComplementForm[24:0]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FADD.scala 129:29]
  wire  result_sign = a_LessThan_b ? ~io_in_a_sign : io_in_a_sign; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FADD.scala 132:24]
  wire [7:0] resultExpNoRound = lza_io_zero ? 8'h0 : io_in_a_exp; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FADD.scala 146:29]
  wire  resultExpIsZero = resultExpNoRound == 8'h0; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FADD.scala 147:42]
  wire [4:0] _GEN_0 = {{4'd0}, lza_io_error}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FADD.scala 149:45]
  wire [4:0] _shiftLimit_T_1 = lza_io_lzc + _GEN_0; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FADD.scala 149:45]
  wire [7:0] _GEN_1 = {{3'd0}, _shiftLimit_T_1}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FADD.scala 149:37]
  wire  shiftLimit = resultExpNoRound <= _GEN_1; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FADD.scala 149:37]
  wire [7:0] _GEN_2 = {{3'd0}, lza_io_lzc}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FADD.scala 150:33]
  wire [7:0] exp_s1 = resultExpNoRound - _GEN_2; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FADD.scala 150:33]
  wire [7:0] _GEN_3 = {{7'd0}, lza_io_error}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FADD.scala 151:23]
  wire [7:0] exp_s2 = exp_s1 - _GEN_3; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FADD.scala 151:23]
  wire [7:0] closePathResult_exp = shiftLimit ? 8'h0 : exp_s2; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FADD.scala 152:29]
  wire [7:0] _sigShiftNum_T_1 = resultExpNoRound - 8'h1; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FADD.scala 157:39]
  wire [7:0] _sigShiftNum_T_2 = shiftLimit ? _sigShiftNum_T_1 : {{3'd0}, lza_io_lzc}; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [7:0] sigShiftNum = resultExpIsZero ? 8'h0 : _sigShiftNum_T_2; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [279:0] _GEN_5 = {{255'd0}, resultSigNoRound}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FADD.scala 161:34]
  wire [279:0] _sig_s1_T = _GEN_5 << sigShiftNum; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FADD.scala 161:34]
  wire [24:0] sig_s1 = _sig_s1_T[24:0]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FADD.scala 161:49]
  wire [24:0] _sig_s2_T_1 = {sig_s1[23:0],1'h0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FADD.scala 162:33]
  wire [24:0] sig_s2 = lza_io_error ? _sig_s2_T_1 : sig_s1; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FADD.scala 162:19]
  wire [24:0] _sig_s3_T = shiftLimit ? sig_s1 : sig_s2; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FADD.scala 165:10]
  wire [26:0] sig_s3 = {_sig_s3_T,2'h0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FADD.scala 164:8]
  wire [26:0] close_path_sig = {sig_s3[26:1],|sig_s3[0]}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FADD.scala 171:53]
  wire [7:0] _GEN_4 = {{7'd0}, near_path_rounder_io_cout}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FADD.scala 186:57]
  wire [7:0] near_path_exp_rounded = _GEN_4 + closePathResult_exp; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FADD.scala 186:57]
  wire  _io_out_result_T_1 = result_sign & ~lza_io_zero; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FADD.scala 190:27]
  wire [8:0] io_out_result_hi = {_io_out_result_T_1,near_path_exp_rounded}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FADD.scala 189:23]
  LZA lza ( // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FADD.scala 134:19]
    .io_a(lza_io_a),
    .io_b(lza_io_b),
    .io_lzc(lza_io_lzc),
    .io_error(lza_io_error),
    .io_zero(lza_io_zero)
  );
  TininessRounder near_path_tininess_rounder ( // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FADD.scala 174:42]
    .io_in_sig(near_path_tininess_rounder_io_in_sig)
  );
  RoundingUnit near_path_rounder ( // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/RoundingUnit.scala 44:25]
    .io_in(near_path_rounder_io_in),
    .io_roundIn(near_path_rounder_io_roundIn),
    .io_stickyIn(near_path_rounder_io_stickyIn),
    .io_out(near_path_rounder_io_out),
    .io_cout(near_path_rounder_io_cout)
  );
  assign io_out_result = {io_out_result_hi,near_path_rounder_io_out}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FADD.scala 189:23]
  assign io_out_near_path_of = near_path_exp_rounded == 8'hff; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FADD.scala 195:48]
  assign lza_io_a = {io_in_a_sig,1'h0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FADD.scala 122:18]
  assign lza_io_b = _b_sig_T >> io_in_needShift; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FADD.scala 123:43]
  assign near_path_tininess_rounder_io_in_sig = {sig_s3[26:1],|sig_s3[0]}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FADD.scala 171:53]
  assign near_path_rounder_io_in = close_path_sig[25:3]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/RoundingUnit.scala 45:33]
  assign near_path_rounder_io_roundIn = close_path_sig[2]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/RoundingUnit.scala 46:50]
  assign near_path_rounder_io_stickyIn = |close_path_sig[1:0]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/RoundingUnit.scala 47:51]
endmodule
module FADD(
  output        io_in_ready, // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FADD.scala 221:14]
  input         io_in_valid, // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FADD.scala 221:14]
  input  [31:0] io_in_bits_a, // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FADD.scala 221:14]
  input  [31:0] io_in_bits_b, // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FADD.scala 221:14]
  input         io_in_bits_a_inter_valid, // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FADD.scala 221:14]
  input         io_in_bits_b_inter_valid, // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FADD.scala 221:14]
  input         io_in_bits_a_inter_flags_isNaN, // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FADD.scala 221:14]
  input         io_in_bits_a_inter_flags_isInf, // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FADD.scala 221:14]
  input         io_in_bits_b_inter_flags_isNaN, // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FADD.scala 221:14]
  input         io_in_bits_b_inter_flags_isInf, // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FADD.scala 221:14]
  input         io_out_ready, // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FADD.scala 221:14]
  output        io_out_valid, // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FADD.scala 221:14]
  output [31:0] io_out_bits_result // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FADD.scala 221:14]
);
  wire  farPath_io_in_a_sign; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FADD.scala 247:23]
  wire [7:0] farPath_io_in_a_exp; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FADD.scala 247:23]
  wire [23:0] farPath_io_in_a_sig; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FADD.scala 247:23]
  wire [7:0] farPath_io_in_b_exp; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FADD.scala 247:23]
  wire [23:0] farPath_io_in_b_sig; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FADD.scala 247:23]
  wire  farPath_io_in_addSig; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FADD.scala 247:23]
  wire  farPath_io_in_tinyAdd; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FADD.scala 247:23]
  wire [4:0] farPath_io_in_shiftNum; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FADD.scala 247:23]
  wire [31:0] farPath_io_out_result; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FADD.scala 247:23]
  wire  farPath_io_out_far_path_of; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FADD.scala 247:23]
  wire  closePath_io_in_a_sign; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FADD.scala 261:25]
  wire [7:0] closePath_io_in_a_exp; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FADD.scala 261:25]
  wire [23:0] closePath_io_in_a_sig; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FADD.scala 261:25]
  wire [7:0] closePath_io_in_b_exp; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FADD.scala 261:25]
  wire [23:0] closePath_io_in_b_sig; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FADD.scala 261:25]
  wire  closePath_io_in_needShift; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FADD.scala 261:25]
  wire [31:0] closePath_io_out_result; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FADD.scala 261:25]
  wire  closePath_io_out_near_path_of; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FADD.scala 261:25]
  wire  fp_a_sign = io_in_bits_a[31]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/package.scala 58:19]
  wire [7:0] fp_a_exp = io_in_bits_a[30:23]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/package.scala 59:18]
  wire [22:0] fp_a_sig = io_in_bits_a[22:0]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/package.scala 60:18]
  wire  fp_b_sign = io_in_bits_b[31]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/package.scala 58:19]
  wire [7:0] fp_b_exp = io_in_bits_b[30:23]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/package.scala 59:18]
  wire [22:0] fp_b_sig = io_in_bits_b[22:0]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/package.scala 60:18]
  wire  decode_a_expNotZero = |fp_a_exp; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/package.scala 31:28]
  wire  decode_a_expIsOnes = &fp_a_exp; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/package.scala 32:27]
  wire  decode_a_sigNotZero = |fp_a_sig; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/package.scala 33:28]
  wire  decode_a__expIsZero = ~decode_a_expNotZero; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/package.scala 36:27]
  wire  decode_a__sigIsZero = ~decode_a_sigNotZero; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/package.scala 39:27]
  wire  decode_a__isSubnormal = decode_a__expIsZero & decode_a_sigNotZero; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/package.scala 40:46]
  wire  decode_a__isInf = decode_a_expIsOnes & decode_a__sigIsZero; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/package.scala 41:40]
  wire  decode_a__isNaN = decode_a_expIsOnes & decode_a_sigNotZero; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/package.scala 43:40]
  wire  decode_b_expNotZero = |fp_b_exp; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/package.scala 31:28]
  wire  decode_b_expIsOnes = &fp_b_exp; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/package.scala 32:27]
  wire  decode_b_sigNotZero = |fp_b_sig; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/package.scala 33:28]
  wire  decode_b__expIsZero = ~decode_b_expNotZero; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/package.scala 36:27]
  wire  decode_b__sigIsZero = ~decode_b_sigNotZero; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/package.scala 39:27]
  wire  decode_b__isSubnormal = decode_b__expIsZero & decode_b_sigNotZero; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/package.scala 40:46]
  wire  decode_b__isInf = decode_b_expIsOnes & decode_b__sigIsZero; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/package.scala 41:40]
  wire  decode_b__isNaN = decode_b_expIsOnes & decode_b_sigNotZero; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/package.scala 43:40]
  wire [7:0] _raw_a_inner_exp_T_1 = fp_a_exp + 8'h1; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/package.scala 83:38]
  wire [7:0] raw_a_exp = decode_a__isSubnormal ? _raw_a_inner_exp_T_1 : fp_a_exp; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/package.scala 83:23]
  wire [23:0] raw_a_sig = {decode_a_expNotZero,fp_a_sig}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/package.scala 84:23]
  wire [7:0] _raw_b_inner_exp_T_1 = fp_b_exp + 8'h1; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/package.scala 83:38]
  wire [7:0] raw_b_exp = decode_b__isSubnormal ? _raw_b_inner_exp_T_1 : fp_b_exp; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/package.scala 83:23]
  wire [23:0] raw_b_sig = {decode_b_expNotZero,fp_b_sig}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/package.scala 84:23]
  wire  addSig = fp_a_sign == fp_b_sign; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FADD.scala 235:26]
  wire  needSwap = raw_a_exp < raw_b_exp; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FADD.scala 236:28]
  wire [7:0] _diffExp_T_1 = raw_b_exp - raw_a_exp; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FADD.scala 237:41]
  wire [7:0] _diffExp_T_3 = raw_a_exp - raw_b_exp; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FADD.scala 237:64]
  wire [7:0] diffExp = needSwap ? _diffExp_T_1 : _diffExp_T_3; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FADD.scala 237:20]
  wire [4:0] initShiftNum = diffExp[4:0]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FADD.scala 240:29]
  wire  isMaxAlign = diffExp > 8'h1a; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FADD.scala 241:28]
  wire  _closePathSel_T = ~addSig; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FADD.scala 243:22]
  wire  closePathSel = ~addSig & ~isMaxAlign & initShiftNum <= 5'h1; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FADD.scala 243:45]
  wire  a_isNaN = io_in_bits_a_inter_valid ? io_in_bits_a_inter_flags_isNaN : decode_a__isNaN; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FADD.scala 275:20]
  wire  a_isInf = io_in_bits_a_inter_valid ? io_in_bits_a_inter_flags_isInf : decode_a__isInf; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FADD.scala 277:20]
  wire  b_isNaN = io_in_bits_b_inter_valid ? io_in_bits_b_inter_flags_isNaN : decode_b__isNaN; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FADD.scala 281:20]
  wire  b_isInf = io_in_bits_b_inter_valid ? io_in_bits_b_inter_flags_isInf : decode_b__isInf; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FADD.scala 283:20]
  wire  special_path_hasNaN = a_isNaN | b_isNaN; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FADD.scala 285:37]
  wire  special_path_hasInf = a_isInf | b_isInf; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FADD.scala 287:37]
  wire  special_path_inf_iv = a_isInf & b_isInf & _closePathSel_T; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FADD.scala 288:48]
  wire  special_case_happen = special_path_hasNaN | special_path_hasInf; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FADD.scala 289:49]
  wire  _special_path_result_T = special_path_hasNaN | special_path_inf_iv; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FADD.scala 293:25]
  wire  _special_path_result_T_3 = a_isInf ? fp_a_sign : fp_b_sign; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FADD.scala 296:10]
  wire [31:0] _special_path_result_T_5 = {_special_path_result_T_3,8'hff,23'h0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FADD.scala 295:8]
  wire [31:0] special_path_result = _special_path_result_T ? 32'h7fc00000 : _special_path_result_T_5; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FADD.scala 292:32]
  wire  common_overflow_sign = closePathSel ? closePath_io_out_result[31] : farPath_io_out_result[31]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FADD.scala 306:8]
  wire  common_overflow = ~closePathSel & farPath_io_out_far_path_of | closePathSel & closePath_io_out_near_path_of; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FADD.scala 316:34]
  wire [31:0] _io_out_bits_result_T = {common_overflow_sign,8'hff,23'h0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FADD.scala 336:10]
  wire [31:0] _io_out_bits_result_T_1 = closePathSel ? closePath_io_out_result : farPath_io_out_result; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FADD.scala 337:10]
  wire [31:0] _io_out_bits_result_T_2 = common_overflow ? _io_out_bits_result_T : _io_out_bits_result_T_1; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FADD.scala 334:8]
  FarPath farPath ( // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FADD.scala 247:23]
    .io_in_a_sign(farPath_io_in_a_sign),
    .io_in_a_exp(farPath_io_in_a_exp),
    .io_in_a_sig(farPath_io_in_a_sig),
    .io_in_b_exp(farPath_io_in_b_exp),
    .io_in_b_sig(farPath_io_in_b_sig),
    .io_in_addSig(farPath_io_in_addSig),
    .io_in_tinyAdd(farPath_io_in_tinyAdd),
    .io_in_shiftNum(farPath_io_in_shiftNum),
    .io_out_result(farPath_io_out_result),
    .io_out_far_path_of(farPath_io_out_far_path_of)
  );
  ClosePath closePath ( // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FADD.scala 261:25]
    .io_in_a_sign(closePath_io_in_a_sign),
    .io_in_a_exp(closePath_io_in_a_exp),
    .io_in_a_sig(closePath_io_in_a_sig),
    .io_in_b_exp(closePath_io_in_b_exp),
    .io_in_b_sig(closePath_io_in_b_sig),
    .io_in_needShift(closePath_io_in_needShift),
    .io_out_result(closePath_io_out_result),
    .io_out_near_path_of(closePath_io_out_near_path_of)
  );
  assign io_in_ready = io_out_ready; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FADD.scala 329:15]
  assign io_out_valid = io_in_valid; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FADD.scala 330:16]
  assign io_out_bits_result = special_case_happen ? special_path_result : _io_out_bits_result_T_2; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FADD.scala 331:28]
  assign farPath_io_in_a_sign = needSwap ? fp_b_sign : fp_a_sign; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FADD.scala 248:25]
  assign farPath_io_in_a_exp = needSwap ? raw_b_exp : raw_a_exp; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FADD.scala 248:25]
  assign farPath_io_in_a_sig = needSwap ? raw_b_sig : raw_a_sig; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FADD.scala 248:25]
  assign farPath_io_in_b_exp = needSwap ? raw_a_exp : raw_b_exp; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FADD.scala 249:25]
  assign farPath_io_in_b_sig = needSwap ? raw_a_sig : raw_b_sig; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FADD.scala 249:25]
  assign farPath_io_in_addSig = fp_a_sign == fp_b_sign; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FADD.scala 235:26]
  assign farPath_io_in_tinyAdd = decode_a__expIsZero & decode_b__expIsZero; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FADD.scala 251:47]
  assign farPath_io_in_shiftNum = isMaxAlign ? 5'h1a : initShiftNum; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FADD.scala 242:21]
  assign closePath_io_in_a_sign = needSwap ? fp_b_sign : fp_a_sign; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FADD.scala 262:27]
  assign closePath_io_in_a_exp = needSwap ? raw_b_exp : raw_a_exp; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FADD.scala 262:27]
  assign closePath_io_in_a_sig = needSwap ? raw_b_sig : raw_a_sig; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FADD.scala 262:27]
  assign closePath_io_in_b_exp = needSwap ? raw_a_exp : raw_b_exp; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FADD.scala 263:27]
  assign closePath_io_in_b_sig = needSwap ? raw_a_sig : raw_b_sig; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FADD.scala 263:27]
  assign closePath_io_in_needShift = initShiftNum == 5'h1; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FADD.scala 264:45]
endmodule
module RoundingUnit_16(
  input  [9:0] io_in, // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/RoundingUnit.scala 7:14]
  input        io_roundIn, // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/RoundingUnit.scala 7:14]
  input        io_stickyIn, // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/RoundingUnit.scala 7:14]
  output [9:0] io_out, // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/RoundingUnit.scala 7:14]
  output       io_cout // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/RoundingUnit.scala 7:14]
);
  wire  g = io_in[0]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/RoundingUnit.scala 19:25]
  wire  r_up = io_roundIn & io_stickyIn | io_roundIn & ~io_stickyIn & g; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/RoundingUnit.scala 25:24]
  wire [9:0] out_r_up = io_in + 10'h1; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/RoundingUnit.scala 32:24]
  assign io_out = r_up ? out_r_up : io_in; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/RoundingUnit.scala 33:16]
  assign io_cout = r_up & &io_in; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/RoundingUnit.scala 36:19]
endmodule
module ShiftRightJam_4(
  input  [11:0] io_in, // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/ShiftRightJam.scala 11:14]
  input  [7:0]  io_shamt, // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/ShiftRightJam.scala 11:14]
  output [11:0] io_out, // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/ShiftRightJam.scala 11:14]
  output        io_sticky // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/ShiftRightJam.scala 11:14]
);
  wire  exceed_max_shift = io_shamt > 8'hc; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/ShiftRightJam.scala 17:35]
  wire [3:0] shamt = io_shamt[3:0]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/ShiftRightJam.scala 18:23]
  wire [15:0] _sticky_mask_T = 16'h1 << shamt; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/ShiftRightJam.scala 20:11]
  wire [15:0] _sticky_mask_T_2 = _sticky_mask_T - 16'h1; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/ShiftRightJam.scala 20:28]
  wire [11:0] _sticky_mask_T_5 = exceed_max_shift ? 12'hfff : 12'h0; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/ShiftRightJam.scala 20:53]
  wire [11:0] sticky_mask = _sticky_mask_T_2[11:0] | _sticky_mask_T_5; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/ShiftRightJam.scala 20:47]
  wire [11:0] _io_out_T = io_in >> io_shamt; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/ShiftRightJam.scala 21:46]
  wire [11:0] _io_sticky_T = io_in & sticky_mask; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/ShiftRightJam.scala 22:23]
  assign io_out = exceed_max_shift ? 12'h0 : _io_out_T; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/ShiftRightJam.scala 21:16]
  assign io_sticky = |_io_sticky_T; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/ShiftRightJam.scala 22:38]
endmodule
module FPDownConverter(
  input         io_in_valid, // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FPToFP.scala 77:14]
  input  [31:0] io_in_bits_in, // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FPToFP.scala 77:14]
  output        io_out_valid, // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FPToFP.scala 77:14]
  output [15:0] io_out_bits_result // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FPToFP.scala 77:14]
);
  wire [9:0] normal_rounder_io_in; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FPToFP.scala 99:30]
  wire  normal_rounder_io_roundIn; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FPToFP.scala 99:30]
  wire  normal_rounder_io_stickyIn; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FPToFP.scala 99:30]
  wire [9:0] normal_rounder_io_out; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FPToFP.scala 99:30]
  wire  normal_rounder_io_cout; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FPToFP.scala 99:30]
  wire [11:0] shiftRightJam_io_in; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/ShiftRightJam.scala 27:31]
  wire [7:0] shiftRightJam_io_shamt; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/ShiftRightJam.scala 27:31]
  wire [11:0] shiftRightJam_io_out; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/ShiftRightJam.scala 27:31]
  wire  shiftRightJam_io_sticky; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/ShiftRightJam.scala 27:31]
  wire [9:0] subnormal_rounder_io_in; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FPToFP.scala 125:33]
  wire  subnormal_rounder_io_roundIn; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FPToFP.scala 125:33]
  wire  subnormal_rounder_io_stickyIn; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FPToFP.scala 125:33]
  wire [9:0] subnormal_rounder_io_out; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FPToFP.scala 125:33]
  wire  subnormal_rounder_io_cout; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FPToFP.scala 125:33]
  wire  fp_in_sign = io_in_bits_in[31]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/package.scala 58:19]
  wire [7:0] fp_in_exp = io_in_bits_in[30:23]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/package.scala 59:18]
  wire [22:0] fp_in_sig = io_in_bits_in[22:0]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/package.scala 60:18]
  wire  decode_expNotZero = |fp_in_exp; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/package.scala 31:28]
  wire  decode_expIsOnes = &fp_in_exp; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/package.scala 32:27]
  wire  decode_sigNotZero = |fp_in_sig; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/package.scala 33:28]
  wire  decode__isNaN = decode_expIsOnes & decode_sigNotZero; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/package.scala 43:40]
  wire [8:0] _resultExpNoRound_T = {1'b0,$signed(fp_in_exp)}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FPToFP.scala 90:36]
  wire [8:0] resultExpNoRound = $signed(_resultExpNoRound_T) - 9'sh70; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FPToFP.scala 90:41]
  wire  normal_stickyBit = |fp_in_sig[11:0]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FPToFP.scala 97:54]
  wire [8:0] _normal_exp_rounded_T_2 = $signed(resultExpNoRound) + 9'sh1; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FPToFP.scala 107:73]
  wire [8:0] normal_exp_rounded = normal_rounder_io_cout ? $signed(_normal_exp_rounded_T_2) : $signed(resultExpNoRound); // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FPToFP.scala 107:31]
  wire  _expOverflow_T = $signed(resultExpNoRound) > 9'sh1d; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FPToFP.scala 110:22]
  wire  _expOverflow_T_1 = $signed(resultExpNoRound) > 9'sh1e; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FPToFP.scala 111:22]
  wire  expOverflow = normal_rounder_io_cout ? _expOverflow_T : _expOverflow_T_1; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FPToFP.scala 108:24]
  wire  _expUnderflow_T_1 = $signed(resultExpNoRound) < 9'sh1; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FPToFP.scala 113:91]
  wire  subnormal_exp_rounded = subnormal_rounder_io_cout; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FPToFP.scala 132:34]
  wire  _common_exp_T = ~_expUnderflow_T_1; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FPToFP.scala 153:7]
  wire  _common_exp_T_1 = ~_expUnderflow_T_1 & expOverflow; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FPToFP.scala 153:23]
  wire  _common_exp_T_4 = _common_exp_T & ~expOverflow; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FPToFP.scala 154:23]
  wire [4:0] _common_exp_T_6 = _common_exp_T_1 ? 5'h1f : 5'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [4:0] _common_exp_T_7 = _common_exp_T_4 ? normal_exp_rounded[4:0] : 5'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _common_exp_T_8 = _expUnderflow_T_1 & subnormal_exp_rounded; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [4:0] _common_exp_T_9 = _common_exp_T_6 | _common_exp_T_7; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [4:0] _GEN_0 = {{4'd0}, _common_exp_T_8}; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [4:0] common_exp = _common_exp_T_9 | _GEN_0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [9:0] _common_sig_T_6 = _common_exp_T_4 ? normal_rounder_io_out : 10'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [9:0] _common_sig_T_7 = _expUnderflow_T_1 ? subnormal_rounder_io_out : 10'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [9:0] common_sig = _common_sig_T_6 | _common_sig_T_7; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _of_T = ~decode_expIsOnes; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FPToFP.scala 182:12]
  wire  _result_T_1 = ~decode__isNaN & fp_in_sign; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FPToFP.scala 192:19]
  wire [4:0] _result_T_4 = decode_expIsOnes ? 5'h1f : 5'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [4:0] _result_T_5 = _of_T ? common_exp : 5'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [4:0] _result_T_6 = _result_T_4 | _result_T_5; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [9:0] _result_T_8 = {decode_sigNotZero,9'h0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FPToFP.scala 200:12]
  wire [9:0] _result_T_9 = decode_expIsOnes ? _result_T_8 : 10'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [9:0] _result_T_10 = _of_T ? common_sig : 10'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [9:0] _result_T_11 = _result_T_9 | _result_T_10; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [5:0] result_hi = {_result_T_1,_result_T_6}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FPToFP.scala 191:19]
  RoundingUnit_16 normal_rounder ( // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FPToFP.scala 99:30]
    .io_in(normal_rounder_io_in),
    .io_roundIn(normal_rounder_io_roundIn),
    .io_stickyIn(normal_rounder_io_stickyIn),
    .io_out(normal_rounder_io_out),
    .io_cout(normal_rounder_io_cout)
  );
  ShiftRightJam_4 shiftRightJam ( // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/ShiftRightJam.scala 27:31]
    .io_in(shiftRightJam_io_in),
    .io_shamt(shiftRightJam_io_shamt),
    .io_out(shiftRightJam_io_out),
    .io_sticky(shiftRightJam_io_sticky)
  );
  RoundingUnit_16 subnormal_rounder ( // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FPToFP.scala 125:33]
    .io_in(subnormal_rounder_io_in),
    .io_roundIn(subnormal_rounder_io_roundIn),
    .io_stickyIn(subnormal_rounder_io_stickyIn),
    .io_out(subnormal_rounder_io_out),
    .io_cout(subnormal_rounder_io_cout)
  );
  assign io_out_valid = io_in_valid; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FPToFP.scala 207:16]
  assign io_out_bits_result = {result_hi,_result_T_11}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FPToFP.scala 191:19]
  assign normal_rounder_io_in = fp_in_sig[22:13]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FPToFP.scala 95:34]
  assign normal_rounder_io_roundIn = fp_in_sig[12]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FPToFP.scala 96:61]
  assign normal_rounder_io_stickyIn = |fp_in_sig[11:0]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FPToFP.scala 97:54]
  assign shiftRightJam_io_in = {decode_expNotZero,fp_in_sig[22:12]}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FPToFP.scala 121:8]
  assign shiftRightJam_io_shamt = 8'h71 - fp_in_exp; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FPToFP.scala 119:45]
  assign subnormal_rounder_io_in = shiftRightJam_io_out[10:1]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FPToFP.scala 126:56]
  assign subnormal_rounder_io_roundIn = shiftRightJam_io_out[0]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FPToFP.scala 127:48]
  assign subnormal_rounder_io_stickyIn = shiftRightJam_io_sticky | normal_stickyBit; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FPToFP.scala 124:42]
endmodule
module DotProdUnit(
  input         clock,
  input         reset,
  output        io_in_ready, // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/DotProdUnit.scala 30:14]
  input         io_in_valid, // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/DotProdUnit.scala 30:14]
  input  [15:0] io_in_bits_vec_a_0, // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/DotProdUnit.scala 30:14]
  input  [15:0] io_in_bits_vec_a_1, // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/DotProdUnit.scala 30:14]
  input  [15:0] io_in_bits_vec_a_2, // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/DotProdUnit.scala 30:14]
  input  [15:0] io_in_bits_vec_a_3, // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/DotProdUnit.scala 30:14]
  input  [15:0] io_in_bits_vec_b_0, // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/DotProdUnit.scala 30:14]
  input  [15:0] io_in_bits_vec_b_1, // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/DotProdUnit.scala 30:14]
  input  [15:0] io_in_bits_vec_b_2, // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/DotProdUnit.scala 30:14]
  input  [15:0] io_in_bits_vec_b_3, // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/DotProdUnit.scala 30:14]
  input  [31:0] io_in_bits_c, // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/DotProdUnit.scala 30:14]
  input         io_in_bits_mixPc, // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/DotProdUnit.scala 30:14]
  input  [1:0]  io_in_bits_rowtag, // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/DotProdUnit.scala 30:14]
  output        io_out_valid, // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/DotProdUnit.scala 30:14]
  output [31:0] io_out_bits_result, // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/DotProdUnit.scala 30:14]
  output        io_out_bits_mixPc, // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/DotProdUnit.scala 30:14]
  output [1:0]  io_out_bits_rowtag // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/DotProdUnit.scala 30:14]
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
`endif // RANDOMIZE_REG_INIT
  wire  fmul_io_in_ready; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FMUL.scala 106:22]
  wire  fmul_io_in_valid; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FMUL.scala 106:22]
  wire [15:0] fmul_io_in_bits_a; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FMUL.scala 106:22]
  wire [15:0] fmul_io_in_bits_b; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FMUL.scala 106:22]
  wire  fmul_io_toFADD_ready; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FMUL.scala 106:22]
  wire  fmul_io_toFADD_valid; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FMUL.scala 106:22]
  wire [31:0] fmul_io_toFADD_bits_fp_prod; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FMUL.scala 106:22]
  wire  fmul_io_toFADD_bits_inter_flags_isNaN; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FMUL.scala 106:22]
  wire  fmul_io_toFADD_bits_inter_flags_isInf; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FMUL.scala 106:22]
  wire  fmul_1_io_in_ready; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FMUL.scala 106:22]
  wire  fmul_1_io_in_valid; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FMUL.scala 106:22]
  wire [15:0] fmul_1_io_in_bits_a; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FMUL.scala 106:22]
  wire [15:0] fmul_1_io_in_bits_b; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FMUL.scala 106:22]
  wire  fmul_1_io_toFADD_ready; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FMUL.scala 106:22]
  wire  fmul_1_io_toFADD_valid; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FMUL.scala 106:22]
  wire [31:0] fmul_1_io_toFADD_bits_fp_prod; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FMUL.scala 106:22]
  wire  fmul_1_io_toFADD_bits_inter_flags_isNaN; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FMUL.scala 106:22]
  wire  fmul_1_io_toFADD_bits_inter_flags_isInf; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FMUL.scala 106:22]
  wire  fmul_2_io_in_ready; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FMUL.scala 106:22]
  wire  fmul_2_io_in_valid; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FMUL.scala 106:22]
  wire [15:0] fmul_2_io_in_bits_a; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FMUL.scala 106:22]
  wire [15:0] fmul_2_io_in_bits_b; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FMUL.scala 106:22]
  wire  fmul_2_io_toFADD_ready; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FMUL.scala 106:22]
  wire  fmul_2_io_toFADD_valid; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FMUL.scala 106:22]
  wire [31:0] fmul_2_io_toFADD_bits_fp_prod; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FMUL.scala 106:22]
  wire  fmul_2_io_toFADD_bits_inter_flags_isNaN; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FMUL.scala 106:22]
  wire  fmul_2_io_toFADD_bits_inter_flags_isInf; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FMUL.scala 106:22]
  wire  fmul_3_io_in_ready; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FMUL.scala 106:22]
  wire  fmul_3_io_in_valid; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FMUL.scala 106:22]
  wire [15:0] fmul_3_io_in_bits_a; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FMUL.scala 106:22]
  wire [15:0] fmul_3_io_in_bits_b; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FMUL.scala 106:22]
  wire  fmul_3_io_toFADD_ready; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FMUL.scala 106:22]
  wire  fmul_3_io_toFADD_valid; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FMUL.scala 106:22]
  wire [31:0] fmul_3_io_toFADD_bits_fp_prod; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FMUL.scala 106:22]
  wire  fmul_3_io_toFADD_bits_inter_flags_isNaN; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FMUL.scala 106:22]
  wire  fmul_3_io_toFADD_bits_inter_flags_isInf; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FMUL.scala 106:22]
  wire  fcvt_io_in_ready; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FPToFP.scala 314:22]
  wire [15:0] fcvt_io_in_bits_in; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FPToFP.scala 314:22]
  wire  fcvt_io_out_ready; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FPToFP.scala 314:22]
  wire [31:0] fcvt_io_out_bits_result; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FPToFP.scala 314:22]
  wire  faddModule_io_in_ready; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FADD.scala 352:28]
  wire  faddModule_io_in_valid; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FADD.scala 352:28]
  wire [31:0] faddModule_io_in_bits_a; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FADD.scala 352:28]
  wire [31:0] faddModule_io_in_bits_b; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FADD.scala 352:28]
  wire  faddModule_io_in_bits_a_inter_valid; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FADD.scala 352:28]
  wire  faddModule_io_in_bits_b_inter_valid; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FADD.scala 352:28]
  wire  faddModule_io_in_bits_a_inter_flags_isNaN; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FADD.scala 352:28]
  wire  faddModule_io_in_bits_a_inter_flags_isInf; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FADD.scala 352:28]
  wire  faddModule_io_in_bits_b_inter_flags_isNaN; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FADD.scala 352:28]
  wire  faddModule_io_in_bits_b_inter_flags_isInf; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FADD.scala 352:28]
  wire  faddModule_io_out_ready; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FADD.scala 352:28]
  wire  faddModule_io_out_valid; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FADD.scala 352:28]
  wire [31:0] faddModule_io_out_bits_result; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FADD.scala 352:28]
  wire  faddModule_1_io_in_ready; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FADD.scala 352:28]
  wire  faddModule_1_io_in_valid; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FADD.scala 352:28]
  wire [31:0] faddModule_1_io_in_bits_a; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FADD.scala 352:28]
  wire [31:0] faddModule_1_io_in_bits_b; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FADD.scala 352:28]
  wire  faddModule_1_io_in_bits_a_inter_valid; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FADD.scala 352:28]
  wire  faddModule_1_io_in_bits_b_inter_valid; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FADD.scala 352:28]
  wire  faddModule_1_io_in_bits_a_inter_flags_isNaN; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FADD.scala 352:28]
  wire  faddModule_1_io_in_bits_a_inter_flags_isInf; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FADD.scala 352:28]
  wire  faddModule_1_io_in_bits_b_inter_flags_isNaN; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FADD.scala 352:28]
  wire  faddModule_1_io_in_bits_b_inter_flags_isInf; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FADD.scala 352:28]
  wire  faddModule_1_io_out_ready; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FADD.scala 352:28]
  wire  faddModule_1_io_out_valid; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FADD.scala 352:28]
  wire [31:0] faddModule_1_io_out_bits_result; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FADD.scala 352:28]
  wire  faddModule_2_io_in_ready; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FADD.scala 352:28]
  wire  faddModule_2_io_in_valid; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FADD.scala 352:28]
  wire [31:0] faddModule_2_io_in_bits_a; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FADD.scala 352:28]
  wire [31:0] faddModule_2_io_in_bits_b; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FADD.scala 352:28]
  wire  faddModule_2_io_in_bits_a_inter_valid; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FADD.scala 352:28]
  wire  faddModule_2_io_in_bits_b_inter_valid; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FADD.scala 352:28]
  wire  faddModule_2_io_in_bits_a_inter_flags_isNaN; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FADD.scala 352:28]
  wire  faddModule_2_io_in_bits_a_inter_flags_isInf; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FADD.scala 352:28]
  wire  faddModule_2_io_in_bits_b_inter_flags_isNaN; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FADD.scala 352:28]
  wire  faddModule_2_io_in_bits_b_inter_flags_isInf; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FADD.scala 352:28]
  wire  faddModule_2_io_out_ready; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FADD.scala 352:28]
  wire  faddModule_2_io_out_valid; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FADD.scala 352:28]
  wire [31:0] faddModule_2_io_out_bits_result; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FADD.scala 352:28]
  wire  faddModule_3_io_in_ready; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FADD.scala 352:28]
  wire  faddModule_3_io_in_valid; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FADD.scala 352:28]
  wire [31:0] faddModule_3_io_in_bits_a; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FADD.scala 352:28]
  wire [31:0] faddModule_3_io_in_bits_b; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FADD.scala 352:28]
  wire  faddModule_3_io_in_bits_a_inter_valid; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FADD.scala 352:28]
  wire  faddModule_3_io_in_bits_b_inter_valid; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FADD.scala 352:28]
  wire  faddModule_3_io_in_bits_a_inter_flags_isNaN; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FADD.scala 352:28]
  wire  faddModule_3_io_in_bits_a_inter_flags_isInf; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FADD.scala 352:28]
  wire  faddModule_3_io_in_bits_b_inter_flags_isNaN; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FADD.scala 352:28]
  wire  faddModule_3_io_in_bits_b_inter_flags_isInf; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FADD.scala 352:28]
  wire  faddModule_3_io_out_ready; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FADD.scala 352:28]
  wire  faddModule_3_io_out_valid; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FADD.scala 352:28]
  wire [31:0] faddModule_3_io_out_bits_result; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FADD.scala 352:28]
  wire  fcvt_1_io_in_valid; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FPToFP.scala 220:22]
  wire [31:0] fcvt_1_io_in_bits_in; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FPToFP.scala 220:22]
  wire  fcvt_1_io_out_valid; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FPToFP.scala 220:22]
  wire [15:0] fcvt_1_io_out_bits_result; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FPToFP.scala 220:22]
  wire  firstFaddReady_0 = faddModule_io_in_ready; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/DotProdUnit.scala 49:28 85:25]
  wire  firstFaddReady_1 = faddModule_1_io_in_ready; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/DotProdUnit.scala 49:28 85:25]
  wire  _T = firstFaddReady_0 & firstFaddReady_1; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/DotProdUnit.scala 51:134]
  wire  fmulReady_0 = fmul_io_in_ready; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/DotProdUnit.scala 46:34 54:18]
  wire  fmulReady_1 = fmul_1_io_in_ready; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/DotProdUnit.scala 46:34 54:18]
  wire  fmulReady_2 = fmul_2_io_in_ready; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/DotProdUnit.scala 46:34 54:18]
  wire  fmulReady_3 = fmul_3_io_in_ready; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/DotProdUnit.scala 46:34 54:18]
  wire  fmulValid_0 = fmul_io_toFADD_valid; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/DotProdUnit.scala 46:34 53:18]
  wire  fmulValid_1 = fmul_1_io_toFADD_valid; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/DotProdUnit.scala 46:34 53:18]
  wire  _s1_handshaked_s2_T = fmulValid_0 & fmulValid_1; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/DotProdUnit.scala 66:44]
  wire  fmulValid_2 = fmul_2_io_toFADD_valid; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/DotProdUnit.scala 46:34 53:18]
  wire  fmulValid_3 = fmul_3_io_toFADD_valid; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/DotProdUnit.scala 46:34 53:18]
  wire  s1_handshaked_s2 = fmulValid_0 & fmulValid_1 & fmulValid_2 & fmulValid_3 & _T; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/DotProdUnit.scala 66:49]
  reg  mixPc_s2; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/DotProdUnit.scala 67:27]
  reg [1:0] rowtag_s2; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/DotProdUnit.scala 69:28]
  wire  prehandshaked = _s1_handshaked_s2_T & faddModule_io_in_ready; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FADD.scala 354:35]
  reg  valid; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FADD.scala 355:24]
  wire  firstPostReady_0 = faddModule_2_io_in_ready; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/DotProdUnit.scala 117:23 72:28]
  wire  _GEN_3 = faddModule_io_out_valid & firstPostReady_0 ? 1'h0 : valid; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FADD.scala 356:49 357:13 355:24]
  wire  _GEN_4 = prehandshaked | _GEN_3; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FADD.scala 359:25 360:13]
  reg  a_flag_isNaN; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FADD.scala 365:55]
  reg  a_flag_isInf; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FADD.scala 365:55]
  wire  fmulResult_0_inter_flags_isNaN = fmul_io_toFADD_bits_inter_flags_isNaN; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/DotProdUnit.scala 45:24 52:19]
  wire  fmulResult_0_inter_flags_isInf = fmul_io_toFADD_bits_inter_flags_isInf; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/DotProdUnit.scala 45:24 52:19]
  reg  b_flag_isNaN; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FADD.scala 366:55]
  reg  b_flag_isInf; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FADD.scala 366:55]
  wire  fmulResult_1_inter_flags_isNaN = fmul_1_io_toFADD_bits_inter_flags_isNaN; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/DotProdUnit.scala 45:24 52:19]
  wire  fmulResult_1_inter_flags_isInf = fmul_1_io_toFADD_bits_inter_flags_isInf; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/DotProdUnit.scala 45:24 52:19]
  reg [31:0] faddModule_io_in_bits_a_r; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FADD.scala 370:41]
  wire [31:0] fmulResult_0_fp_prod = fmul_io_toFADD_bits_fp_prod; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/DotProdUnit.scala 45:24 52:19]
  reg [31:0] faddModule_io_in_bits_b_r; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FADD.scala 371:41]
  wire [31:0] fmulResult_1_fp_prod = fmul_1_io_toFADD_bits_fp_prod; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/DotProdUnit.scala 45:24 52:19]
  wire  prevalid_1 = fmulValid_2 & fmulValid_3; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/DotProdUnit.scala 79:39]
  wire  prehandshaked_1 = prevalid_1 & faddModule_1_io_in_ready; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FADD.scala 354:35]
  reg  valid_1; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FADD.scala 355:24]
  wire  _GEN_15 = faddModule_1_io_out_valid & firstPostReady_0 ? 1'h0 : valid_1; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FADD.scala 356:49 357:13 355:24]
  wire  _GEN_16 = prehandshaked_1 | _GEN_15; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FADD.scala 359:25 360:13]
  reg  a_flag_1_isNaN; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FADD.scala 365:55]
  reg  a_flag_1_isInf; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FADD.scala 365:55]
  wire  fmulResult_2_inter_flags_isNaN = fmul_2_io_toFADD_bits_inter_flags_isNaN; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/DotProdUnit.scala 45:24 52:19]
  wire  fmulResult_2_inter_flags_isInf = fmul_2_io_toFADD_bits_inter_flags_isInf; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/DotProdUnit.scala 45:24 52:19]
  reg  b_flag_1_isNaN; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FADD.scala 366:55]
  reg  b_flag_1_isInf; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FADD.scala 366:55]
  wire  fmulResult_3_inter_flags_isNaN = fmul_3_io_toFADD_bits_inter_flags_isNaN; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/DotProdUnit.scala 45:24 52:19]
  wire  fmulResult_3_inter_flags_isInf = fmul_3_io_toFADD_bits_inter_flags_isInf; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/DotProdUnit.scala 45:24 52:19]
  reg [31:0] faddModule_io_in_bits_a_r_1; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FADD.scala 370:41]
  wire [31:0] fmulResult_2_fp_prod = fmul_2_io_toFADD_bits_fp_prod; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/DotProdUnit.scala 45:24 52:19]
  reg [31:0] faddModule_io_in_bits_b_r_1; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FADD.scala 371:41]
  wire [31:0] fmulResult_3_fp_prod = fmul_3_io_toFADD_bits_fp_prod; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/DotProdUnit.scala 45:24 52:19]
  reg [31:0] firstAddResult_2_r; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/DotProdUnit.scala 90:45]
  wire  firstFaddValid_0 = faddModule_io_out_valid; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/DotProdUnit.scala 71:28 84:25]
  wire  firstFaddValid_1 = faddModule_1_io_out_valid; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/DotProdUnit.scala 71:28 84:25]
  wire  _T_13 = firstFaddValid_0 & firstFaddValid_1; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/DotProdUnit.scala 134:124]
  wire  prehandshaked_2 = _T_13 & firstPostReady_0; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/DotProdUnit.scala 96:34]
  reg  mixPc_this; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/DotProdUnit.scala 98:31]
  reg [1:0] rowtag_this; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/DotProdUnit.scala 99:32]
  wire  prehandshaked_3 = _T_13 & faddModule_2_io_in_ready; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FADD.scala 354:35]
  reg  valid_2; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FADD.scala 355:24]
  wire  postReady_0 = faddModule_3_io_in_ready; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/DotProdUnit.scala 109:27 128:22]
  wire  _GEN_31 = faddModule_2_io_out_valid & postReady_0 ? 1'h0 : valid_2; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FADD.scala 356:49 357:13 355:24]
  wire  _GEN_32 = prehandshaked_3 | _GEN_31; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FADD.scala 359:25 360:13]
  reg [31:0] faddModule_io_in_bits_a_r_2; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FADD.scala 370:41]
  wire [31:0] firstAddResult_0 = faddModule_io_out_bits_result; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/DotProdUnit.scala 70:28 83:25]
  reg [31:0] faddModule_io_in_bits_b_r_2; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FADD.scala 371:41]
  wire [31:0] firstAddResult_1 = faddModule_1_io_out_bits_result; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/DotProdUnit.scala 70:28 83:25]
  reg [31:0] addResult_1_r; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/DotProdUnit.scala 119:36]
  wire  postValid_0 = faddModule_2_io_out_valid; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/DotProdUnit.scala 108:27 116:24]
  wire  posthandshaked = postValid_0 & postReady_0; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/DotProdUnit.scala 123:53]
  reg  mixPc_sx; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/DotProdUnit.scala 125:36]
  reg [1:0] rowtag_sx; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/DotProdUnit.scala 126:37]
  wire  prehandshaked_4 = postValid_0 & faddModule_3_io_in_ready; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FADD.scala 354:35]
  reg  valid_3; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FADD.scala 355:24]
  wire  _T_15 = faddModule_3_io_out_valid; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FADD.scala 356:34]
  wire  _GEN_39 = faddModule_3_io_out_valid ? 1'h0 : valid_3; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FADD.scala 356:49 357:13 355:24]
  wire  _GEN_40 = prehandshaked_4 | _GEN_39; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FADD.scala 359:25 360:13]
  reg [31:0] faddModule_io_in_bits_a_r_3; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FADD.scala 370:41]
  wire [31:0] addResult_0 = faddModule_2_io_out_bits_result; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/DotProdUnit.scala 107:27 115:24]
  reg [31:0] faddModule_io_in_bits_b_r_3; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FADD.scala 371:41]
  reg  mixPc_es; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/DotProdUnit.scala 141:27]
  reg [1:0] rowtag_es; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/DotProdUnit.scala 142:28]
  reg [31:0] atResult_es; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/DotProdUnit.scala 143:30]
  reg  esValid; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/DotProdUnit.scala 146:24]
  wire  _GEN_48 = io_out_valid ? 1'h0 : esValid; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/DotProdUnit.scala 147:22 148:13 146:24]
  wire  _GEN_49 = _T_15 | _GEN_48; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/DotProdUnit.scala 150:25 151:13]
  wire  prehandshaked_5 = faddModule_3_io_out_valid & ~mixPc_sx; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/DotProdUnit.scala 154:110]
  reg  valid_4; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FPToFP.scala 223:24]
  wire  _GEN_50 = fcvt_1_io_out_valid ? 1'h0 : valid_4; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FPToFP.scala 224:43 225:13 223:24]
  wire  _GEN_51 = prehandshaked_5 | _GEN_50; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FPToFP.scala 227:25 228:13]
  reg [31:0] fcvt_io_in_bits_in_r; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FPToFP.scala 232:36]
  wire [15:0] _io_out_bits_result_T_1 = fcvt_1_io_out_bits_result; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/package.scala 94:22]
  wire [31:0] _io_out_bits_result_T_2 = {16'hffff,_io_out_bits_result_T_1}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/package.scala 94:8]
  FMULnoRound fmul ( // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FMUL.scala 106:22]
    .io_in_ready(fmul_io_in_ready),
    .io_in_valid(fmul_io_in_valid),
    .io_in_bits_a(fmul_io_in_bits_a),
    .io_in_bits_b(fmul_io_in_bits_b),
    .io_toFADD_ready(fmul_io_toFADD_ready),
    .io_toFADD_valid(fmul_io_toFADD_valid),
    .io_toFADD_bits_fp_prod(fmul_io_toFADD_bits_fp_prod),
    .io_toFADD_bits_inter_flags_isNaN(fmul_io_toFADD_bits_inter_flags_isNaN),
    .io_toFADD_bits_inter_flags_isInf(fmul_io_toFADD_bits_inter_flags_isInf)
  );
  FMULnoRound fmul_1 ( // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FMUL.scala 106:22]
    .io_in_ready(fmul_1_io_in_ready),
    .io_in_valid(fmul_1_io_in_valid),
    .io_in_bits_a(fmul_1_io_in_bits_a),
    .io_in_bits_b(fmul_1_io_in_bits_b),
    .io_toFADD_ready(fmul_1_io_toFADD_ready),
    .io_toFADD_valid(fmul_1_io_toFADD_valid),
    .io_toFADD_bits_fp_prod(fmul_1_io_toFADD_bits_fp_prod),
    .io_toFADD_bits_inter_flags_isNaN(fmul_1_io_toFADD_bits_inter_flags_isNaN),
    .io_toFADD_bits_inter_flags_isInf(fmul_1_io_toFADD_bits_inter_flags_isInf)
  );
  FMULnoRound fmul_2 ( // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FMUL.scala 106:22]
    .io_in_ready(fmul_2_io_in_ready),
    .io_in_valid(fmul_2_io_in_valid),
    .io_in_bits_a(fmul_2_io_in_bits_a),
    .io_in_bits_b(fmul_2_io_in_bits_b),
    .io_toFADD_ready(fmul_2_io_toFADD_ready),
    .io_toFADD_valid(fmul_2_io_toFADD_valid),
    .io_toFADD_bits_fp_prod(fmul_2_io_toFADD_bits_fp_prod),
    .io_toFADD_bits_inter_flags_isNaN(fmul_2_io_toFADD_bits_inter_flags_isNaN),
    .io_toFADD_bits_inter_flags_isInf(fmul_2_io_toFADD_bits_inter_flags_isInf)
  );
  FMULnoRound fmul_3 ( // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FMUL.scala 106:22]
    .io_in_ready(fmul_3_io_in_ready),
    .io_in_valid(fmul_3_io_in_valid),
    .io_in_bits_a(fmul_3_io_in_bits_a),
    .io_in_bits_b(fmul_3_io_in_bits_b),
    .io_toFADD_ready(fmul_3_io_toFADD_ready),
    .io_toFADD_valid(fmul_3_io_toFADD_valid),
    .io_toFADD_bits_fp_prod(fmul_3_io_toFADD_bits_fp_prod),
    .io_toFADD_bits_inter_flags_isNaN(fmul_3_io_toFADD_bits_inter_flags_isNaN),
    .io_toFADD_bits_inter_flags_isInf(fmul_3_io_toFADD_bits_inter_flags_isInf)
  );
  FPUpConverter fcvt ( // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FPToFP.scala 314:22]
    .io_in_ready(fcvt_io_in_ready),
    .io_in_bits_in(fcvt_io_in_bits_in),
    .io_out_ready(fcvt_io_out_ready),
    .io_out_bits_result(fcvt_io_out_bits_result)
  );
  FADD faddModule ( // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FADD.scala 352:28]
    .io_in_ready(faddModule_io_in_ready),
    .io_in_valid(faddModule_io_in_valid),
    .io_in_bits_a(faddModule_io_in_bits_a),
    .io_in_bits_b(faddModule_io_in_bits_b),
    .io_in_bits_a_inter_valid(faddModule_io_in_bits_a_inter_valid),
    .io_in_bits_b_inter_valid(faddModule_io_in_bits_b_inter_valid),
    .io_in_bits_a_inter_flags_isNaN(faddModule_io_in_bits_a_inter_flags_isNaN),
    .io_in_bits_a_inter_flags_isInf(faddModule_io_in_bits_a_inter_flags_isInf),
    .io_in_bits_b_inter_flags_isNaN(faddModule_io_in_bits_b_inter_flags_isNaN),
    .io_in_bits_b_inter_flags_isInf(faddModule_io_in_bits_b_inter_flags_isInf),
    .io_out_ready(faddModule_io_out_ready),
    .io_out_valid(faddModule_io_out_valid),
    .io_out_bits_result(faddModule_io_out_bits_result)
  );
  FADD faddModule_1 ( // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FADD.scala 352:28]
    .io_in_ready(faddModule_1_io_in_ready),
    .io_in_valid(faddModule_1_io_in_valid),
    .io_in_bits_a(faddModule_1_io_in_bits_a),
    .io_in_bits_b(faddModule_1_io_in_bits_b),
    .io_in_bits_a_inter_valid(faddModule_1_io_in_bits_a_inter_valid),
    .io_in_bits_b_inter_valid(faddModule_1_io_in_bits_b_inter_valid),
    .io_in_bits_a_inter_flags_isNaN(faddModule_1_io_in_bits_a_inter_flags_isNaN),
    .io_in_bits_a_inter_flags_isInf(faddModule_1_io_in_bits_a_inter_flags_isInf),
    .io_in_bits_b_inter_flags_isNaN(faddModule_1_io_in_bits_b_inter_flags_isNaN),
    .io_in_bits_b_inter_flags_isInf(faddModule_1_io_in_bits_b_inter_flags_isInf),
    .io_out_ready(faddModule_1_io_out_ready),
    .io_out_valid(faddModule_1_io_out_valid),
    .io_out_bits_result(faddModule_1_io_out_bits_result)
  );
  FADD faddModule_2 ( // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FADD.scala 352:28]
    .io_in_ready(faddModule_2_io_in_ready),
    .io_in_valid(faddModule_2_io_in_valid),
    .io_in_bits_a(faddModule_2_io_in_bits_a),
    .io_in_bits_b(faddModule_2_io_in_bits_b),
    .io_in_bits_a_inter_valid(faddModule_2_io_in_bits_a_inter_valid),
    .io_in_bits_b_inter_valid(faddModule_2_io_in_bits_b_inter_valid),
    .io_in_bits_a_inter_flags_isNaN(faddModule_2_io_in_bits_a_inter_flags_isNaN),
    .io_in_bits_a_inter_flags_isInf(faddModule_2_io_in_bits_a_inter_flags_isInf),
    .io_in_bits_b_inter_flags_isNaN(faddModule_2_io_in_bits_b_inter_flags_isNaN),
    .io_in_bits_b_inter_flags_isInf(faddModule_2_io_in_bits_b_inter_flags_isInf),
    .io_out_ready(faddModule_2_io_out_ready),
    .io_out_valid(faddModule_2_io_out_valid),
    .io_out_bits_result(faddModule_2_io_out_bits_result)
  );
  FADD faddModule_3 ( // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FADD.scala 352:28]
    .io_in_ready(faddModule_3_io_in_ready),
    .io_in_valid(faddModule_3_io_in_valid),
    .io_in_bits_a(faddModule_3_io_in_bits_a),
    .io_in_bits_b(faddModule_3_io_in_bits_b),
    .io_in_bits_a_inter_valid(faddModule_3_io_in_bits_a_inter_valid),
    .io_in_bits_b_inter_valid(faddModule_3_io_in_bits_b_inter_valid),
    .io_in_bits_a_inter_flags_isNaN(faddModule_3_io_in_bits_a_inter_flags_isNaN),
    .io_in_bits_a_inter_flags_isInf(faddModule_3_io_in_bits_a_inter_flags_isInf),
    .io_in_bits_b_inter_flags_isNaN(faddModule_3_io_in_bits_b_inter_flags_isNaN),
    .io_in_bits_b_inter_flags_isInf(faddModule_3_io_in_bits_b_inter_flags_isInf),
    .io_out_ready(faddModule_3_io_out_ready),
    .io_out_valid(faddModule_3_io_out_valid),
    .io_out_bits_result(faddModule_3_io_out_bits_result)
  );
  FPDownConverter fcvt_1 ( // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FPToFP.scala 220:22]
    .io_in_valid(fcvt_1_io_in_valid),
    .io_in_bits_in(fcvt_1_io_in_bits_in),
    .io_out_valid(fcvt_1_io_out_valid),
    .io_out_bits_result(fcvt_1_io_out_bits_result)
  );
  assign io_in_ready = fmulReady_0 & fmulReady_1 & fmulReady_2 & fmulReady_3 & fcvt_io_in_ready; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/DotProdUnit.scala 62:41]
  assign io_out_valid = fcvt_1_io_out_valid | mixPc_es & esValid; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/DotProdUnit.scala 159:32]
  assign io_out_bits_result = mixPc_es ? atResult_es : _io_out_bits_result_T_2; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/DotProdUnit.scala 155:28]
  assign io_out_bits_mixPc = mixPc_es; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/DotProdUnit.scala 157:21]
  assign io_out_bits_rowtag = rowtag_es; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/DotProdUnit.scala 158:22]
  assign fmul_io_in_valid = io_in_valid; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FMUL.scala 117:22]
  assign fmul_io_in_bits_a = io_in_bits_vec_a_0; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FMUL.scala 120:23]
  assign fmul_io_in_bits_b = io_in_bits_vec_b_0; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FMUL.scala 121:23]
  assign fmul_io_toFADD_ready = firstFaddReady_0 & firstFaddReady_1; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/DotProdUnit.scala 51:134]
  assign fmul_1_io_in_valid = io_in_valid; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FMUL.scala 117:22]
  assign fmul_1_io_in_bits_a = io_in_bits_vec_a_1; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FMUL.scala 120:23]
  assign fmul_1_io_in_bits_b = io_in_bits_vec_b_1; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FMUL.scala 121:23]
  assign fmul_1_io_toFADD_ready = firstFaddReady_0 & firstFaddReady_1; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/DotProdUnit.scala 51:134]
  assign fmul_2_io_in_valid = io_in_valid; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FMUL.scala 117:22]
  assign fmul_2_io_in_bits_a = io_in_bits_vec_a_2; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FMUL.scala 120:23]
  assign fmul_2_io_in_bits_b = io_in_bits_vec_b_2; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FMUL.scala 121:23]
  assign fmul_2_io_toFADD_ready = firstFaddReady_0 & firstFaddReady_1; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/DotProdUnit.scala 51:134]
  assign fmul_3_io_in_valid = io_in_valid; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FMUL.scala 117:22]
  assign fmul_3_io_in_bits_a = io_in_bits_vec_a_3; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FMUL.scala 120:23]
  assign fmul_3_io_in_bits_b = io_in_bits_vec_b_3; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FMUL.scala 121:23]
  assign fmul_3_io_toFADD_ready = firstFaddReady_0 & firstFaddReady_1; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/DotProdUnit.scala 51:134]
  assign fcvt_io_in_bits_in = &io_in_bits_c[31:16] ? io_in_bits_c[15:0] : 16'h7e00; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/package.scala 87:8]
  assign fcvt_io_out_ready = firstFaddReady_0 & firstFaddReady_1; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/DotProdUnit.scala 57:124]
  assign faddModule_io_in_valid = valid; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FADD.scala 368:28]
  assign faddModule_io_in_bits_a = faddModule_io_in_bits_a_r; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FADD.scala 370:29]
  assign faddModule_io_in_bits_b = faddModule_io_in_bits_b_r; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FADD.scala 371:29]
  assign faddModule_io_in_bits_a_inter_valid = 1'h1; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FADD.scala 373:41]
  assign faddModule_io_in_bits_b_inter_valid = 1'h1; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FADD.scala 374:41]
  assign faddModule_io_in_bits_a_inter_flags_isNaN = a_flag_isNaN; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FADD.scala 375:41]
  assign faddModule_io_in_bits_a_inter_flags_isInf = a_flag_isInf; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FADD.scala 375:41]
  assign faddModule_io_in_bits_b_inter_flags_isNaN = b_flag_isNaN; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FADD.scala 376:41]
  assign faddModule_io_in_bits_b_inter_flags_isInf = b_flag_isInf; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FADD.scala 376:41]
  assign faddModule_io_out_ready = faddModule_2_io_in_ready; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/DotProdUnit.scala 117:23 72:28]
  assign faddModule_1_io_in_valid = valid_1; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FADD.scala 368:28]
  assign faddModule_1_io_in_bits_a = faddModule_io_in_bits_a_r_1; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FADD.scala 370:29]
  assign faddModule_1_io_in_bits_b = faddModule_io_in_bits_b_r_1; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FADD.scala 371:29]
  assign faddModule_1_io_in_bits_a_inter_valid = 1'h1; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FADD.scala 373:41]
  assign faddModule_1_io_in_bits_b_inter_valid = 1'h1; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FADD.scala 374:41]
  assign faddModule_1_io_in_bits_a_inter_flags_isNaN = a_flag_1_isNaN; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FADD.scala 375:41]
  assign faddModule_1_io_in_bits_a_inter_flags_isInf = a_flag_1_isInf; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FADD.scala 375:41]
  assign faddModule_1_io_in_bits_b_inter_flags_isNaN = b_flag_1_isNaN; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FADD.scala 376:41]
  assign faddModule_1_io_in_bits_b_inter_flags_isInf = b_flag_1_isInf; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FADD.scala 376:41]
  assign faddModule_1_io_out_ready = faddModule_2_io_in_ready; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/DotProdUnit.scala 117:23 72:28]
  assign faddModule_2_io_in_valid = valid_2; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FADD.scala 368:28]
  assign faddModule_2_io_in_bits_a = faddModule_io_in_bits_a_r_2; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FADD.scala 370:29]
  assign faddModule_2_io_in_bits_b = faddModule_io_in_bits_b_r_2; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FADD.scala 371:29]
  assign faddModule_2_io_in_bits_a_inter_valid = 1'h0; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FADD.scala 373:41]
  assign faddModule_2_io_in_bits_b_inter_valid = 1'h0; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FADD.scala 374:41]
  assign faddModule_2_io_in_bits_a_inter_flags_isNaN = 1'h0;
  assign faddModule_2_io_in_bits_a_inter_flags_isInf = 1'h0;
  assign faddModule_2_io_in_bits_b_inter_flags_isNaN = 1'h0;
  assign faddModule_2_io_in_bits_b_inter_flags_isInf = 1'h0;
  assign faddModule_2_io_out_ready = faddModule_3_io_in_ready; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/DotProdUnit.scala 109:27 128:22]
  assign faddModule_3_io_in_valid = valid_3; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FADD.scala 368:28]
  assign faddModule_3_io_in_bits_a = faddModule_io_in_bits_a_r_3; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FADD.scala 370:29]
  assign faddModule_3_io_in_bits_b = faddModule_io_in_bits_b_r_3; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FADD.scala 371:29]
  assign faddModule_3_io_in_bits_a_inter_valid = 1'h0; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FADD.scala 373:41]
  assign faddModule_3_io_in_bits_b_inter_valid = 1'h0; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FADD.scala 374:41]
  assign faddModule_3_io_in_bits_a_inter_flags_isNaN = 1'h0;
  assign faddModule_3_io_in_bits_a_inter_flags_isInf = 1'h0;
  assign faddModule_3_io_in_bits_b_inter_flags_isNaN = 1'h0;
  assign faddModule_3_io_in_bits_b_inter_flags_isInf = 1'h0;
  assign faddModule_3_io_out_ready = 1'h1; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FADD.scala 377:29]
  assign fcvt_1_io_in_valid = valid_4; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FPToFP.scala 231:22]
  assign fcvt_1_io_in_bits_in = fcvt_io_in_bits_in_r; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FPToFP.scala 232:24]
  always @(posedge clock) begin
    if (s1_handshaked_s2) begin // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/DotProdUnit.scala 67:27]
      mixPc_s2 <= io_in_bits_mixPc; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/DotProdUnit.scala 67:27]
    end
    if (s1_handshaked_s2) begin // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/DotProdUnit.scala 69:28]
      rowtag_s2 <= io_in_bits_rowtag; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/DotProdUnit.scala 69:28]
    end
    if (reset) begin // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FADD.scala 355:24]
      valid <= 1'h0; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FADD.scala 355:24]
    end else begin
      valid <= _GEN_4;
    end
    if (prehandshaked) begin // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FADD.scala 365:55]
      a_flag_isNaN <= fmulResult_0_inter_flags_isNaN; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FADD.scala 365:55]
    end
    if (prehandshaked) begin // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FADD.scala 365:55]
      a_flag_isInf <= fmulResult_0_inter_flags_isInf; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FADD.scala 365:55]
    end
    if (prehandshaked) begin // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FADD.scala 366:55]
      b_flag_isNaN <= fmulResult_1_inter_flags_isNaN; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FADD.scala 366:55]
    end
    if (prehandshaked) begin // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FADD.scala 366:55]
      b_flag_isInf <= fmulResult_1_inter_flags_isInf; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FADD.scala 366:55]
    end
    if (prehandshaked) begin // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FADD.scala 370:41]
      faddModule_io_in_bits_a_r <= fmulResult_0_fp_prod; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FADD.scala 370:41]
    end
    if (prehandshaked) begin // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FADD.scala 371:41]
      faddModule_io_in_bits_b_r <= fmulResult_1_fp_prod; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FADD.scala 371:41]
    end
    if (reset) begin // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FADD.scala 355:24]
      valid_1 <= 1'h0; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FADD.scala 355:24]
    end else begin
      valid_1 <= _GEN_16;
    end
    if (prehandshaked_1) begin // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FADD.scala 365:55]
      a_flag_1_isNaN <= fmulResult_2_inter_flags_isNaN; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FADD.scala 365:55]
    end
    if (prehandshaked_1) begin // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FADD.scala 365:55]
      a_flag_1_isInf <= fmulResult_2_inter_flags_isInf; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FADD.scala 365:55]
    end
    if (prehandshaked_1) begin // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FADD.scala 366:55]
      b_flag_1_isNaN <= fmulResult_3_inter_flags_isNaN; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FADD.scala 366:55]
    end
    if (prehandshaked_1) begin // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FADD.scala 366:55]
      b_flag_1_isInf <= fmulResult_3_inter_flags_isInf; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FADD.scala 366:55]
    end
    if (prehandshaked_1) begin // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FADD.scala 370:41]
      faddModule_io_in_bits_a_r_1 <= fmulResult_2_fp_prod; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FADD.scala 370:41]
    end
    if (prehandshaked_1) begin // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FADD.scala 371:41]
      faddModule_io_in_bits_b_r_1 <= fmulResult_3_fp_prod; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FADD.scala 371:41]
    end
    if (s1_handshaked_s2) begin // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/DotProdUnit.scala 90:45]
      if (io_in_bits_mixPc) begin // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/DotProdUnit.scala 58:19]
        firstAddResult_2_r <= io_in_bits_c;
      end else begin
        firstAddResult_2_r <= fcvt_io_out_bits_result;
      end
    end
    if (prehandshaked_2) begin // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/DotProdUnit.scala 98:31]
      mixPc_this <= mixPc_s2; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/DotProdUnit.scala 98:31]
    end
    if (prehandshaked_2) begin // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/DotProdUnit.scala 99:32]
      rowtag_this <= rowtag_s2; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/DotProdUnit.scala 99:32]
    end
    if (reset) begin // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FADD.scala 355:24]
      valid_2 <= 1'h0; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FADD.scala 355:24]
    end else begin
      valid_2 <= _GEN_32;
    end
    if (prehandshaked_3) begin // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FADD.scala 370:41]
      faddModule_io_in_bits_a_r_2 <= firstAddResult_0; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FADD.scala 370:41]
    end
    if (prehandshaked_3) begin // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FADD.scala 371:41]
      faddModule_io_in_bits_b_r_2 <= firstAddResult_1; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FADD.scala 371:41]
    end
    if (prehandshaked_2) begin // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/DotProdUnit.scala 119:36]
      addResult_1_r <= firstAddResult_2_r; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/DotProdUnit.scala 119:36]
    end
    if (posthandshaked) begin // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/DotProdUnit.scala 125:36]
      mixPc_sx <= mixPc_this; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/DotProdUnit.scala 125:36]
    end
    if (posthandshaked) begin // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/DotProdUnit.scala 126:37]
      rowtag_sx <= rowtag_this; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/DotProdUnit.scala 126:37]
    end
    if (reset) begin // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FADD.scala 355:24]
      valid_3 <= 1'h0; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FADD.scala 355:24]
    end else begin
      valid_3 <= _GEN_40;
    end
    if (prehandshaked_4) begin // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FADD.scala 370:41]
      faddModule_io_in_bits_a_r_3 <= addResult_0; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FADD.scala 370:41]
    end
    if (prehandshaked_4) begin // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FADD.scala 371:41]
      faddModule_io_in_bits_b_r_3 <= addResult_1_r; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FADD.scala 371:41]
    end
    if (_T_15) begin // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/DotProdUnit.scala 141:27]
      mixPc_es <= mixPc_sx; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/DotProdUnit.scala 141:27]
    end
    if (_T_15) begin // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/DotProdUnit.scala 142:28]
      rowtag_es <= rowtag_sx; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/DotProdUnit.scala 142:28]
    end
    if (_T_15) begin // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/DotProdUnit.scala 143:30]
      atResult_es <= faddModule_3_io_out_bits_result; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/DotProdUnit.scala 143:30]
    end
    if (reset) begin // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/DotProdUnit.scala 146:24]
      esValid <= 1'h0; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/DotProdUnit.scala 146:24]
    end else begin
      esValid <= _GEN_49;
    end
    if (reset) begin // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FPToFP.scala 223:24]
      valid_4 <= 1'h0; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FPToFP.scala 223:24]
    end else begin
      valid_4 <= _GEN_51;
    end
    if (prehandshaked_5) begin // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FPToFP.scala 232:36]
      fcvt_io_in_bits_in_r <= faddModule_3_io_out_bits_result; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/fpu/FPToFP.scala 232:36]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  mixPc_s2 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  rowtag_s2 = _RAND_1[1:0];
  _RAND_2 = {1{`RANDOM}};
  valid = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  a_flag_isNaN = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  a_flag_isInf = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  b_flag_isNaN = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  b_flag_isInf = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  faddModule_io_in_bits_a_r = _RAND_7[31:0];
  _RAND_8 = {1{`RANDOM}};
  faddModule_io_in_bits_b_r = _RAND_8[31:0];
  _RAND_9 = {1{`RANDOM}};
  valid_1 = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  a_flag_1_isNaN = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  a_flag_1_isInf = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  b_flag_1_isNaN = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  b_flag_1_isInf = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  faddModule_io_in_bits_a_r_1 = _RAND_14[31:0];
  _RAND_15 = {1{`RANDOM}};
  faddModule_io_in_bits_b_r_1 = _RAND_15[31:0];
  _RAND_16 = {1{`RANDOM}};
  firstAddResult_2_r = _RAND_16[31:0];
  _RAND_17 = {1{`RANDOM}};
  mixPc_this = _RAND_17[0:0];
  _RAND_18 = {1{`RANDOM}};
  rowtag_this = _RAND_18[1:0];
  _RAND_19 = {1{`RANDOM}};
  valid_2 = _RAND_19[0:0];
  _RAND_20 = {1{`RANDOM}};
  faddModule_io_in_bits_a_r_2 = _RAND_20[31:0];
  _RAND_21 = {1{`RANDOM}};
  faddModule_io_in_bits_b_r_2 = _RAND_21[31:0];
  _RAND_22 = {1{`RANDOM}};
  addResult_1_r = _RAND_22[31:0];
  _RAND_23 = {1{`RANDOM}};
  mixPc_sx = _RAND_23[0:0];
  _RAND_24 = {1{`RANDOM}};
  rowtag_sx = _RAND_24[1:0];
  _RAND_25 = {1{`RANDOM}};
  valid_3 = _RAND_25[0:0];
  _RAND_26 = {1{`RANDOM}};
  faddModule_io_in_bits_a_r_3 = _RAND_26[31:0];
  _RAND_27 = {1{`RANDOM}};
  faddModule_io_in_bits_b_r_3 = _RAND_27[31:0];
  _RAND_28 = {1{`RANDOM}};
  mixPc_es = _RAND_28[0:0];
  _RAND_29 = {1{`RANDOM}};
  rowtag_es = _RAND_29[1:0];
  _RAND_30 = {1{`RANDOM}};
  atResult_es = _RAND_30[31:0];
  _RAND_31 = {1{`RANDOM}};
  esValid = _RAND_31[0:0];
  _RAND_32 = {1{`RANDOM}};
  valid_4 = _RAND_32[0:0];
  _RAND_33 = {1{`RANDOM}};
  fcvt_io_in_bits_in_r = _RAND_33[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Threadgroup(
  input          clock,
  input          reset,
  output         io_in_ready, // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/Threadgroup.scala 20:14]
  input          io_in_valid, // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/Threadgroup.scala 20:14]
  input  [255:0] io_in_bits_matrix_a_data, // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/Threadgroup.scala 20:14]
  input  [255:0] io_in_bits_matrix_b_data, // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/Threadgroup.scala 20:14]
  input  [255:0] io_in_bits_matrix_c_data, // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/Threadgroup.scala 20:14]
  input          io_in_bits_mixPcMode, // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/Threadgroup.scala 20:14]
  output         io_out_valid, // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/Threadgroup.scala 20:14]
  output [255:0] io_out_bits_matrix_d_data // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/Threadgroup.scala 20:14]
);
`ifdef RANDOMIZE_REG_INIT
  reg [63:0] _RAND_0;
  reg [63:0] _RAND_1;
  reg [63:0] _RAND_2;
  reg [63:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
`endif // RANDOMIZE_REG_INIT
  wire  dp_clock; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/DotProdUnit.scala 167:20]
  wire  dp_reset; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/DotProdUnit.scala 167:20]
  wire  dp_io_in_ready; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/DotProdUnit.scala 167:20]
  wire  dp_io_in_valid; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/DotProdUnit.scala 167:20]
  wire [15:0] dp_io_in_bits_vec_a_0; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/DotProdUnit.scala 167:20]
  wire [15:0] dp_io_in_bits_vec_a_1; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/DotProdUnit.scala 167:20]
  wire [15:0] dp_io_in_bits_vec_a_2; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/DotProdUnit.scala 167:20]
  wire [15:0] dp_io_in_bits_vec_a_3; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/DotProdUnit.scala 167:20]
  wire [15:0] dp_io_in_bits_vec_b_0; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/DotProdUnit.scala 167:20]
  wire [15:0] dp_io_in_bits_vec_b_1; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/DotProdUnit.scala 167:20]
  wire [15:0] dp_io_in_bits_vec_b_2; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/DotProdUnit.scala 167:20]
  wire [15:0] dp_io_in_bits_vec_b_3; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/DotProdUnit.scala 167:20]
  wire [31:0] dp_io_in_bits_c; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/DotProdUnit.scala 167:20]
  wire  dp_io_in_bits_mixPc; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/DotProdUnit.scala 167:20]
  wire [1:0] dp_io_in_bits_rowtag; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/DotProdUnit.scala 167:20]
  wire  dp_io_out_valid; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/DotProdUnit.scala 167:20]
  wire [31:0] dp_io_out_bits_result; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/DotProdUnit.scala 167:20]
  wire  dp_io_out_bits_mixPc; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/DotProdUnit.scala 167:20]
  wire [1:0] dp_io_out_bits_rowtag; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/DotProdUnit.scala 167:20]
  wire  dp_1_clock; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/DotProdUnit.scala 167:20]
  wire  dp_1_reset; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/DotProdUnit.scala 167:20]
  wire  dp_1_io_in_ready; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/DotProdUnit.scala 167:20]
  wire  dp_1_io_in_valid; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/DotProdUnit.scala 167:20]
  wire [15:0] dp_1_io_in_bits_vec_a_0; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/DotProdUnit.scala 167:20]
  wire [15:0] dp_1_io_in_bits_vec_a_1; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/DotProdUnit.scala 167:20]
  wire [15:0] dp_1_io_in_bits_vec_a_2; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/DotProdUnit.scala 167:20]
  wire [15:0] dp_1_io_in_bits_vec_a_3; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/DotProdUnit.scala 167:20]
  wire [15:0] dp_1_io_in_bits_vec_b_0; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/DotProdUnit.scala 167:20]
  wire [15:0] dp_1_io_in_bits_vec_b_1; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/DotProdUnit.scala 167:20]
  wire [15:0] dp_1_io_in_bits_vec_b_2; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/DotProdUnit.scala 167:20]
  wire [15:0] dp_1_io_in_bits_vec_b_3; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/DotProdUnit.scala 167:20]
  wire [31:0] dp_1_io_in_bits_c; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/DotProdUnit.scala 167:20]
  wire  dp_1_io_in_bits_mixPc; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/DotProdUnit.scala 167:20]
  wire [1:0] dp_1_io_in_bits_rowtag; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/DotProdUnit.scala 167:20]
  wire  dp_1_io_out_valid; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/DotProdUnit.scala 167:20]
  wire [31:0] dp_1_io_out_bits_result; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/DotProdUnit.scala 167:20]
  wire  dp_1_io_out_bits_mixPc; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/DotProdUnit.scala 167:20]
  wire [1:0] dp_1_io_out_bits_rowtag; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/DotProdUnit.scala 167:20]
  wire  dp_2_clock; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/DotProdUnit.scala 167:20]
  wire  dp_2_reset; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/DotProdUnit.scala 167:20]
  wire  dp_2_io_in_ready; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/DotProdUnit.scala 167:20]
  wire  dp_2_io_in_valid; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/DotProdUnit.scala 167:20]
  wire [15:0] dp_2_io_in_bits_vec_a_0; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/DotProdUnit.scala 167:20]
  wire [15:0] dp_2_io_in_bits_vec_a_1; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/DotProdUnit.scala 167:20]
  wire [15:0] dp_2_io_in_bits_vec_a_2; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/DotProdUnit.scala 167:20]
  wire [15:0] dp_2_io_in_bits_vec_a_3; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/DotProdUnit.scala 167:20]
  wire [15:0] dp_2_io_in_bits_vec_b_0; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/DotProdUnit.scala 167:20]
  wire [15:0] dp_2_io_in_bits_vec_b_1; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/DotProdUnit.scala 167:20]
  wire [15:0] dp_2_io_in_bits_vec_b_2; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/DotProdUnit.scala 167:20]
  wire [15:0] dp_2_io_in_bits_vec_b_3; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/DotProdUnit.scala 167:20]
  wire [31:0] dp_2_io_in_bits_c; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/DotProdUnit.scala 167:20]
  wire  dp_2_io_in_bits_mixPc; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/DotProdUnit.scala 167:20]
  wire [1:0] dp_2_io_in_bits_rowtag; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/DotProdUnit.scala 167:20]
  wire  dp_2_io_out_valid; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/DotProdUnit.scala 167:20]
  wire [31:0] dp_2_io_out_bits_result; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/DotProdUnit.scala 167:20]
  wire  dp_2_io_out_bits_mixPc; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/DotProdUnit.scala 167:20]
  wire [1:0] dp_2_io_out_bits_rowtag; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/DotProdUnit.scala 167:20]
  wire  dp_3_clock; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/DotProdUnit.scala 167:20]
  wire  dp_3_reset; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/DotProdUnit.scala 167:20]
  wire  dp_3_io_in_ready; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/DotProdUnit.scala 167:20]
  wire  dp_3_io_in_valid; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/DotProdUnit.scala 167:20]
  wire [15:0] dp_3_io_in_bits_vec_a_0; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/DotProdUnit.scala 167:20]
  wire [15:0] dp_3_io_in_bits_vec_a_1; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/DotProdUnit.scala 167:20]
  wire [15:0] dp_3_io_in_bits_vec_a_2; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/DotProdUnit.scala 167:20]
  wire [15:0] dp_3_io_in_bits_vec_a_3; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/DotProdUnit.scala 167:20]
  wire [15:0] dp_3_io_in_bits_vec_b_0; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/DotProdUnit.scala 167:20]
  wire [15:0] dp_3_io_in_bits_vec_b_1; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/DotProdUnit.scala 167:20]
  wire [15:0] dp_3_io_in_bits_vec_b_2; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/DotProdUnit.scala 167:20]
  wire [15:0] dp_3_io_in_bits_vec_b_3; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/DotProdUnit.scala 167:20]
  wire [31:0] dp_3_io_in_bits_c; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/DotProdUnit.scala 167:20]
  wire  dp_3_io_in_bits_mixPc; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/DotProdUnit.scala 167:20]
  wire [1:0] dp_3_io_in_bits_rowtag; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/DotProdUnit.scala 167:20]
  wire  dp_3_io_out_valid; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/DotProdUnit.scala 167:20]
  wire [31:0] dp_3_io_out_bits_result; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/DotProdUnit.scala 167:20]
  wire  dp_3_io_out_bits_mixPc; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/DotProdUnit.scala 167:20]
  wire [1:0] dp_3_io_out_bits_rowtag; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/DotProdUnit.scala 167:20]
  wire  prehandshaked = io_in_valid & io_in_ready; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/Threadgroup.scala 25:35]
  reg [63:0] matrix_d_0; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/Threadgroup.scala 32:21]
  reg [63:0] matrix_d_1; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/Threadgroup.scala 32:21]
  reg [63:0] matrix_d_2; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/Threadgroup.scala 32:21]
  reg [63:0] matrix_d_3; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/Threadgroup.scala 32:21]
  reg  outValid; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/Threadgroup.scala 38:25]
  wire  _GEN_0 = io_out_valid ? 1'h0 : outValid; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/Threadgroup.scala 39:21 40:14 38:25]
  reg [2:0] state; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/Threadgroup.scala 44:22]
  reg  dp_in_valid; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/Threadgroup.scala 45:28]
  wire [2:0] _GEN_4 = io_in_valid ? 3'h1 : 3'h0; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/Threadgroup.scala 65:33 66:17 68:17]
  wire  _GEN_5 = io_in_valid & dp_in_valid; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/Threadgroup.scala 45:28 65:33 69:23]
  wire [2:0] _GEN_6 = ~io_in_bits_mixPcMode ? 3'h3 : _GEN_4; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/Threadgroup.scala 63:22 64:17]
  wire  _GEN_7 = ~io_in_bits_mixPcMode ? dp_in_valid : _GEN_5; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/Threadgroup.scala 63:22 45:28]
  wire [2:0] _GEN_13 = 3'h4 == state ? _GEN_4 : state; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/Threadgroup.scala 47:17 44:22]
  wire  _GEN_14 = 3'h4 == state ? _GEN_5 : dp_in_valid; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/Threadgroup.scala 47:17 45:28]
  wire [2:0] _GEN_15 = 3'h3 == state ? 3'h4 : _GEN_13; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/Threadgroup.scala 47:17]
  wire  _GEN_16 = 3'h3 == state ? dp_in_valid : _GEN_14; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/Threadgroup.scala 47:17 45:28]
  wire  _dpIn_va_T = state == 3'h2; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/Threadgroup.scala 93:16]
  wire [15:0] dpIn_va_vec__0 = io_in_bits_matrix_a_data[191:176]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/package.scala 44:28]
  wire [15:0] dpIn_va_vec__1 = io_in_bits_matrix_a_data[175:160]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/package.scala 44:28]
  wire [15:0] dpIn_va_vec__2 = io_in_bits_matrix_a_data[159:144]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/package.scala 44:28]
  wire [15:0] dpIn_va_vec__3 = io_in_bits_matrix_a_data[143:128]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/package.scala 44:28]
  wire  _dpIn_va_T_1 = state == 3'h3; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/Threadgroup.scala 94:16]
  wire [15:0] dpIn_va_vec_1_0 = io_in_bits_matrix_a_data[127:112]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/package.scala 44:28]
  wire [15:0] dpIn_va_vec_1_1 = io_in_bits_matrix_a_data[111:96]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/package.scala 44:28]
  wire [15:0] dpIn_va_vec_1_2 = io_in_bits_matrix_a_data[95:80]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/package.scala 44:28]
  wire [15:0] dpIn_va_vec_1_3 = io_in_bits_matrix_a_data[79:64]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/package.scala 44:28]
  wire  _dpIn_va_T_2 = state == 3'h4; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/Threadgroup.scala 95:16]
  wire [15:0] dpIn_va_vec_2_0 = io_in_bits_matrix_a_data[63:48]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/package.scala 44:28]
  wire [15:0] dpIn_va_vec_2_1 = io_in_bits_matrix_a_data[47:32]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/package.scala 44:28]
  wire [15:0] dpIn_va_vec_2_2 = io_in_bits_matrix_a_data[31:16]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/package.scala 44:28]
  wire [15:0] dpIn_va_vec_2_3 = io_in_bits_matrix_a_data[15:0]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/package.scala 44:28]
  wire  _dpIn_va_T_3 = state == 3'h1; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/Threadgroup.scala 96:16]
  wire [15:0] dpIn_va_vec_3_0 = io_in_bits_matrix_a_data[255:240]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/package.scala 44:28]
  wire [15:0] dpIn_va_vec_3_1 = io_in_bits_matrix_a_data[239:224]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/package.scala 44:28]
  wire [15:0] dpIn_va_vec_3_2 = io_in_bits_matrix_a_data[223:208]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/package.scala 44:28]
  wire [15:0] dpIn_va_vec_3_3 = io_in_bits_matrix_a_data[207:192]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/package.scala 44:28]
  wire [15:0] _dpIn_va_T_4 = _dpIn_va_T ? dpIn_va_vec__0 : 16'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [15:0] _dpIn_va_T_5 = _dpIn_va_T_1 ? dpIn_va_vec_1_0 : 16'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [15:0] _dpIn_va_T_6 = _dpIn_va_T_2 ? dpIn_va_vec_2_0 : 16'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [15:0] _dpIn_va_T_7 = _dpIn_va_T_3 ? dpIn_va_vec_3_0 : 16'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [15:0] _dpIn_va_T_8 = _dpIn_va_T_4 | _dpIn_va_T_5; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [15:0] _dpIn_va_T_9 = _dpIn_va_T_8 | _dpIn_va_T_6; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [15:0] _dpIn_va_T_11 = _dpIn_va_T ? dpIn_va_vec__1 : 16'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [15:0] _dpIn_va_T_12 = _dpIn_va_T_1 ? dpIn_va_vec_1_1 : 16'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [15:0] _dpIn_va_T_13 = _dpIn_va_T_2 ? dpIn_va_vec_2_1 : 16'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [15:0] _dpIn_va_T_14 = _dpIn_va_T_3 ? dpIn_va_vec_3_1 : 16'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [15:0] _dpIn_va_T_15 = _dpIn_va_T_11 | _dpIn_va_T_12; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [15:0] _dpIn_va_T_16 = _dpIn_va_T_15 | _dpIn_va_T_13; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [15:0] _dpIn_va_T_18 = _dpIn_va_T ? dpIn_va_vec__2 : 16'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [15:0] _dpIn_va_T_19 = _dpIn_va_T_1 ? dpIn_va_vec_1_2 : 16'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [15:0] _dpIn_va_T_20 = _dpIn_va_T_2 ? dpIn_va_vec_2_2 : 16'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [15:0] _dpIn_va_T_21 = _dpIn_va_T_3 ? dpIn_va_vec_3_2 : 16'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [15:0] _dpIn_va_T_22 = _dpIn_va_T_18 | _dpIn_va_T_19; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [15:0] _dpIn_va_T_23 = _dpIn_va_T_22 | _dpIn_va_T_20; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [15:0] _dpIn_va_T_25 = _dpIn_va_T ? dpIn_va_vec__3 : 16'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [15:0] _dpIn_va_T_26 = _dpIn_va_T_1 ? dpIn_va_vec_1_3 : 16'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [15:0] _dpIn_va_T_27 = _dpIn_va_T_2 ? dpIn_va_vec_2_3 : 16'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [15:0] _dpIn_va_T_28 = _dpIn_va_T_3 ? dpIn_va_vec_3_3 : 16'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [15:0] _dpIn_va_T_29 = _dpIn_va_T_25 | _dpIn_va_T_26; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [15:0] _dpIn_va_T_30 = _dpIn_va_T_29 | _dpIn_va_T_27; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [31:0] dpIn_c_vec__0 = io_in_bits_matrix_c_data[127:96]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/package.scala 44:28]
  wire [31:0] dpIn_c_vec__1 = io_in_bits_matrix_c_data[95:64]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/package.scala 44:28]
  wire [31:0] dpIn_c_vec__2 = io_in_bits_matrix_c_data[63:32]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/package.scala 44:28]
  wire [31:0] dpIn_c_vec__3 = io_in_bits_matrix_c_data[31:0]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/package.scala 44:28]
  wire [15:0] dpIn_c_vec_1_0 = io_in_bits_matrix_c_data[191:176]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/package.scala 44:28]
  wire [15:0] dpIn_c_vec_1_1 = io_in_bits_matrix_c_data[175:160]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/package.scala 44:28]
  wire [15:0] dpIn_c_vec_1_2 = io_in_bits_matrix_c_data[159:144]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/package.scala 44:28]
  wire [15:0] dpIn_c_vec_1_3 = io_in_bits_matrix_c_data[143:128]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/package.scala 44:28]
  wire [31:0] dpIn_c_res_boxed__0 = {16'hffff,dpIn_c_vec_1_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/package.scala 99:26]
  wire [31:0] dpIn_c_res_boxed__1 = {16'hffff,dpIn_c_vec_1_1}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/package.scala 99:26]
  wire [31:0] dpIn_c_res_boxed__2 = {16'hffff,dpIn_c_vec_1_2}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/package.scala 99:26]
  wire [31:0] dpIn_c_res_boxed__3 = {16'hffff,dpIn_c_vec_1_3}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/package.scala 99:26]
  wire [31:0] _dpIn_c_T_1_0 = io_in_bits_mixPcMode ? dpIn_c_vec__0 : dpIn_c_res_boxed__0; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/Threadgroup.scala 102:30]
  wire [31:0] _dpIn_c_T_1_1 = io_in_bits_mixPcMode ? dpIn_c_vec__1 : dpIn_c_res_boxed__1; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/Threadgroup.scala 102:30]
  wire [31:0] _dpIn_c_T_1_2 = io_in_bits_mixPcMode ? dpIn_c_vec__2 : dpIn_c_res_boxed__2; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/Threadgroup.scala 102:30]
  wire [31:0] _dpIn_c_T_1_3 = io_in_bits_mixPcMode ? dpIn_c_vec__3 : dpIn_c_res_boxed__3; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/Threadgroup.scala 102:30]
  wire [15:0] dpIn_c_vec_2_0 = io_in_bits_matrix_c_data[127:112]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/package.scala 44:28]
  wire [15:0] dpIn_c_vec_2_1 = io_in_bits_matrix_c_data[111:96]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/package.scala 44:28]
  wire [15:0] dpIn_c_vec_2_2 = io_in_bits_matrix_c_data[95:80]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/package.scala 44:28]
  wire [15:0] dpIn_c_vec_2_3 = io_in_bits_matrix_c_data[79:64]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/package.scala 44:28]
  wire [31:0] dpIn_c_res_boxed_1_0 = {16'hffff,dpIn_c_vec_2_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/package.scala 99:26]
  wire [31:0] dpIn_c_res_boxed_1_1 = {16'hffff,dpIn_c_vec_2_1}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/package.scala 99:26]
  wire [31:0] dpIn_c_res_boxed_1_2 = {16'hffff,dpIn_c_vec_2_2}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/package.scala 99:26]
  wire [31:0] dpIn_c_res_boxed_1_3 = {16'hffff,dpIn_c_vec_2_3}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/package.scala 99:26]
  wire [15:0] dpIn_c_vec_3_0 = io_in_bits_matrix_c_data[63:48]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/package.scala 44:28]
  wire [15:0] dpIn_c_vec_3_1 = io_in_bits_matrix_c_data[47:32]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/package.scala 44:28]
  wire [15:0] dpIn_c_vec_3_2 = io_in_bits_matrix_c_data[31:16]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/package.scala 44:28]
  wire [15:0] dpIn_c_vec_3_3 = io_in_bits_matrix_c_data[15:0]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/package.scala 44:28]
  wire [31:0] dpIn_c_res_boxed_2_0 = {16'hffff,dpIn_c_vec_3_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/package.scala 99:26]
  wire [31:0] dpIn_c_res_boxed_2_1 = {16'hffff,dpIn_c_vec_3_1}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/package.scala 99:26]
  wire [31:0] dpIn_c_res_boxed_2_2 = {16'hffff,dpIn_c_vec_3_2}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/package.scala 99:26]
  wire [31:0] dpIn_c_res_boxed_2_3 = {16'hffff,dpIn_c_vec_3_3}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/package.scala 99:26]
  wire [31:0] dpIn_c_vec_4_0 = io_in_bits_matrix_c_data[255:224]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/package.scala 44:28]
  wire [31:0] dpIn_c_vec_4_1 = io_in_bits_matrix_c_data[223:192]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/package.scala 44:28]
  wire [31:0] dpIn_c_vec_4_2 = io_in_bits_matrix_c_data[191:160]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/package.scala 44:28]
  wire [31:0] dpIn_c_vec_4_3 = io_in_bits_matrix_c_data[159:128]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/package.scala 44:28]
  wire [15:0] dpIn_c_vec_5_0 = io_in_bits_matrix_c_data[255:240]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/package.scala 44:28]
  wire [15:0] dpIn_c_vec_5_1 = io_in_bits_matrix_c_data[239:224]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/package.scala 44:28]
  wire [15:0] dpIn_c_vec_5_2 = io_in_bits_matrix_c_data[223:208]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/package.scala 44:28]
  wire [15:0] dpIn_c_vec_5_3 = io_in_bits_matrix_c_data[207:192]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/package.scala 44:28]
  wire [31:0] dpIn_c_res_boxed_3_0 = {16'hffff,dpIn_c_vec_5_0}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/package.scala 99:26]
  wire [31:0] dpIn_c_res_boxed_3_1 = {16'hffff,dpIn_c_vec_5_1}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/package.scala 99:26]
  wire [31:0] dpIn_c_res_boxed_3_2 = {16'hffff,dpIn_c_vec_5_2}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/package.scala 99:26]
  wire [31:0] dpIn_c_res_boxed_3_3 = {16'hffff,dpIn_c_vec_5_3}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/package.scala 99:26]
  wire [31:0] _dpIn_c_T_5_0 = io_in_bits_mixPcMode ? dpIn_c_vec_4_0 : dpIn_c_res_boxed_3_0; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/Threadgroup.scala 105:30]
  wire [31:0] _dpIn_c_T_5_1 = io_in_bits_mixPcMode ? dpIn_c_vec_4_1 : dpIn_c_res_boxed_3_1; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/Threadgroup.scala 105:30]
  wire [31:0] _dpIn_c_T_5_2 = io_in_bits_mixPcMode ? dpIn_c_vec_4_2 : dpIn_c_res_boxed_3_2; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/Threadgroup.scala 105:30]
  wire [31:0] _dpIn_c_T_5_3 = io_in_bits_mixPcMode ? dpIn_c_vec_4_3 : dpIn_c_res_boxed_3_3; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/Threadgroup.scala 105:30]
  wire [31:0] _dpIn_c_T_6 = _dpIn_va_T ? _dpIn_c_T_1_0 : 32'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [31:0] _dpIn_c_T_7 = _dpIn_va_T_1 ? dpIn_c_res_boxed_1_0 : 32'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [31:0] _dpIn_c_T_8 = _dpIn_va_T_2 ? dpIn_c_res_boxed_2_0 : 32'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [31:0] _dpIn_c_T_9 = _dpIn_va_T_3 ? _dpIn_c_T_5_0 : 32'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [31:0] _dpIn_c_T_10 = _dpIn_c_T_6 | _dpIn_c_T_7; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [31:0] _dpIn_c_T_11 = _dpIn_c_T_10 | _dpIn_c_T_8; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [31:0] _dpIn_c_T_13 = _dpIn_va_T ? _dpIn_c_T_1_1 : 32'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [31:0] _dpIn_c_T_14 = _dpIn_va_T_1 ? dpIn_c_res_boxed_1_1 : 32'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [31:0] _dpIn_c_T_15 = _dpIn_va_T_2 ? dpIn_c_res_boxed_2_1 : 32'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [31:0] _dpIn_c_T_16 = _dpIn_va_T_3 ? _dpIn_c_T_5_1 : 32'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [31:0] _dpIn_c_T_17 = _dpIn_c_T_13 | _dpIn_c_T_14; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [31:0] _dpIn_c_T_18 = _dpIn_c_T_17 | _dpIn_c_T_15; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [31:0] _dpIn_c_T_20 = _dpIn_va_T ? _dpIn_c_T_1_2 : 32'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [31:0] _dpIn_c_T_21 = _dpIn_va_T_1 ? dpIn_c_res_boxed_1_2 : 32'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [31:0] _dpIn_c_T_22 = _dpIn_va_T_2 ? dpIn_c_res_boxed_2_2 : 32'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [31:0] _dpIn_c_T_23 = _dpIn_va_T_3 ? _dpIn_c_T_5_2 : 32'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [31:0] _dpIn_c_T_24 = _dpIn_c_T_20 | _dpIn_c_T_21; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [31:0] _dpIn_c_T_25 = _dpIn_c_T_24 | _dpIn_c_T_22; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [31:0] _dpIn_c_T_27 = _dpIn_va_T ? _dpIn_c_T_1_3 : 32'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [31:0] _dpIn_c_T_28 = _dpIn_va_T_1 ? dpIn_c_res_boxed_1_3 : 32'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [31:0] _dpIn_c_T_29 = _dpIn_va_T_2 ? dpIn_c_res_boxed_2_3 : 32'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [31:0] _dpIn_c_T_30 = _dpIn_va_T_3 ? _dpIn_c_T_5_3 : 32'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [31:0] _dpIn_c_T_31 = _dpIn_c_T_27 | _dpIn_c_T_28; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [31:0] _dpIn_c_T_32 = _dpIn_c_T_31 | _dpIn_c_T_29; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [1:0] _rowtag_in_T_5 = _dpIn_va_T_1 ? 2'h2 : 2'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [1:0] _rowtag_in_T_6 = _dpIn_va_T_2 ? 2'h3 : 2'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [1:0] _GEN_48 = {{1'd0}, _dpIn_va_T}; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [1:0] _rowtag_in_T_8 = _GEN_48 | _rowtag_in_T_5; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [31:0] dpResult_0 = dp_io_out_bits_result; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/Threadgroup.scala 120:17 31:22]
  wire [31:0] dpResult_1 = dp_1_io_out_bits_result; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/Threadgroup.scala 120:17 31:22]
  wire [31:0] dpResult_2 = dp_2_io_out_bits_result; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/Threadgroup.scala 120:17 31:22]
  wire [31:0] dpResult_3 = dp_3_io_out_bits_result; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/Threadgroup.scala 120:17 31:22]
  wire [63:0] result_fp16 = {dpResult_0[15:0],dpResult_1[15:0],dpResult_2[15:0],dpResult_3[15:0]}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/Threadgroup.scala 128:24]
  wire [63:0] result_fp32_hi = {dpResult_0,dpResult_1}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/Threadgroup.scala 129:27]
  wire [63:0] result_fp32_lo = {dpResult_2,dpResult_3}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/Threadgroup.scala 130:27]
  wire  dpValid_0 = dp_io_out_valid; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/Threadgroup.scala 122:16 34:21]
  wire  dpValid_1 = dp_1_io_out_valid; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/Threadgroup.scala 122:16 34:21]
  wire  dpValid_2 = dp_2_io_out_valid; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/Threadgroup.scala 122:16 34:21]
  wire  dpValid_3 = dp_3_io_out_valid; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/Threadgroup.scala 122:16 34:21]
  wire [1:0] rowtag_out = dp_3_io_out_bits_rowtag; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/Threadgroup.scala 124:16 36:24]
  wire  outMixPc = dp_3_io_out_bits_mixPc; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/Threadgroup.scala 125:14 37:22]
  wire  _GEN_27 = outMixPc | _GEN_0; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/Threadgroup.scala 143:24 146:20]
  wire [63:0] _GEN_29 = 2'h3 == rowtag_out ? result_fp16 : matrix_d_3; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/Threadgroup.scala 133:24 155:21 32:21]
  wire  _GEN_30 = 2'h3 == rowtag_out | _GEN_0; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/Threadgroup.scala 133:24 156:18]
  wire  _GEN_33 = 2'h2 == rowtag_out ? _GEN_0 : _GEN_30; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/Threadgroup.scala 133:24]
  wire [127:0] io_out_bits_matrix_d_data_lo = {matrix_d_2,matrix_d_3}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/Threadgroup.scala 161:35]
  wire [127:0] io_out_bits_matrix_d_data_hi = {matrix_d_0,matrix_d_1}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/Threadgroup.scala 161:35]
  wire  dpReady_0 = dp_io_in_ready; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/Threadgroup.scala 123:16 35:21]
  wire  dpReady_1 = dp_1_io_in_ready; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/Threadgroup.scala 123:16 35:21]
  wire  dpReady_2 = dp_2_io_in_ready; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/Threadgroup.scala 123:16 35:21]
  wire  dpReady_3 = dp_3_io_in_ready; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/Threadgroup.scala 123:16 35:21]
  DotProdUnit dp ( // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/DotProdUnit.scala 167:20]
    .clock(dp_clock),
    .reset(dp_reset),
    .io_in_ready(dp_io_in_ready),
    .io_in_valid(dp_io_in_valid),
    .io_in_bits_vec_a_0(dp_io_in_bits_vec_a_0),
    .io_in_bits_vec_a_1(dp_io_in_bits_vec_a_1),
    .io_in_bits_vec_a_2(dp_io_in_bits_vec_a_2),
    .io_in_bits_vec_a_3(dp_io_in_bits_vec_a_3),
    .io_in_bits_vec_b_0(dp_io_in_bits_vec_b_0),
    .io_in_bits_vec_b_1(dp_io_in_bits_vec_b_1),
    .io_in_bits_vec_b_2(dp_io_in_bits_vec_b_2),
    .io_in_bits_vec_b_3(dp_io_in_bits_vec_b_3),
    .io_in_bits_c(dp_io_in_bits_c),
    .io_in_bits_mixPc(dp_io_in_bits_mixPc),
    .io_in_bits_rowtag(dp_io_in_bits_rowtag),
    .io_out_valid(dp_io_out_valid),
    .io_out_bits_result(dp_io_out_bits_result),
    .io_out_bits_mixPc(dp_io_out_bits_mixPc),
    .io_out_bits_rowtag(dp_io_out_bits_rowtag)
  );
  DotProdUnit dp_1 ( // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/DotProdUnit.scala 167:20]
    .clock(dp_1_clock),
    .reset(dp_1_reset),
    .io_in_ready(dp_1_io_in_ready),
    .io_in_valid(dp_1_io_in_valid),
    .io_in_bits_vec_a_0(dp_1_io_in_bits_vec_a_0),
    .io_in_bits_vec_a_1(dp_1_io_in_bits_vec_a_1),
    .io_in_bits_vec_a_2(dp_1_io_in_bits_vec_a_2),
    .io_in_bits_vec_a_3(dp_1_io_in_bits_vec_a_3),
    .io_in_bits_vec_b_0(dp_1_io_in_bits_vec_b_0),
    .io_in_bits_vec_b_1(dp_1_io_in_bits_vec_b_1),
    .io_in_bits_vec_b_2(dp_1_io_in_bits_vec_b_2),
    .io_in_bits_vec_b_3(dp_1_io_in_bits_vec_b_3),
    .io_in_bits_c(dp_1_io_in_bits_c),
    .io_in_bits_mixPc(dp_1_io_in_bits_mixPc),
    .io_in_bits_rowtag(dp_1_io_in_bits_rowtag),
    .io_out_valid(dp_1_io_out_valid),
    .io_out_bits_result(dp_1_io_out_bits_result),
    .io_out_bits_mixPc(dp_1_io_out_bits_mixPc),
    .io_out_bits_rowtag(dp_1_io_out_bits_rowtag)
  );
  DotProdUnit dp_2 ( // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/DotProdUnit.scala 167:20]
    .clock(dp_2_clock),
    .reset(dp_2_reset),
    .io_in_ready(dp_2_io_in_ready),
    .io_in_valid(dp_2_io_in_valid),
    .io_in_bits_vec_a_0(dp_2_io_in_bits_vec_a_0),
    .io_in_bits_vec_a_1(dp_2_io_in_bits_vec_a_1),
    .io_in_bits_vec_a_2(dp_2_io_in_bits_vec_a_2),
    .io_in_bits_vec_a_3(dp_2_io_in_bits_vec_a_3),
    .io_in_bits_vec_b_0(dp_2_io_in_bits_vec_b_0),
    .io_in_bits_vec_b_1(dp_2_io_in_bits_vec_b_1),
    .io_in_bits_vec_b_2(dp_2_io_in_bits_vec_b_2),
    .io_in_bits_vec_b_3(dp_2_io_in_bits_vec_b_3),
    .io_in_bits_c(dp_2_io_in_bits_c),
    .io_in_bits_mixPc(dp_2_io_in_bits_mixPc),
    .io_in_bits_rowtag(dp_2_io_in_bits_rowtag),
    .io_out_valid(dp_2_io_out_valid),
    .io_out_bits_result(dp_2_io_out_bits_result),
    .io_out_bits_mixPc(dp_2_io_out_bits_mixPc),
    .io_out_bits_rowtag(dp_2_io_out_bits_rowtag)
  );
  DotProdUnit dp_3 ( // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/DotProdUnit.scala 167:20]
    .clock(dp_3_clock),
    .reset(dp_3_reset),
    .io_in_ready(dp_3_io_in_ready),
    .io_in_valid(dp_3_io_in_valid),
    .io_in_bits_vec_a_0(dp_3_io_in_bits_vec_a_0),
    .io_in_bits_vec_a_1(dp_3_io_in_bits_vec_a_1),
    .io_in_bits_vec_a_2(dp_3_io_in_bits_vec_a_2),
    .io_in_bits_vec_a_3(dp_3_io_in_bits_vec_a_3),
    .io_in_bits_vec_b_0(dp_3_io_in_bits_vec_b_0),
    .io_in_bits_vec_b_1(dp_3_io_in_bits_vec_b_1),
    .io_in_bits_vec_b_2(dp_3_io_in_bits_vec_b_2),
    .io_in_bits_vec_b_3(dp_3_io_in_bits_vec_b_3),
    .io_in_bits_c(dp_3_io_in_bits_c),
    .io_in_bits_mixPc(dp_3_io_in_bits_mixPc),
    .io_in_bits_rowtag(dp_3_io_in_bits_rowtag),
    .io_out_valid(dp_3_io_out_valid),
    .io_out_bits_result(dp_3_io_out_bits_result),
    .io_out_bits_mixPc(dp_3_io_out_bits_mixPc),
    .io_out_bits_rowtag(dp_3_io_out_bits_rowtag)
  );
  assign io_in_ready = dpReady_0 & dpReady_1 & dpReady_2 & dpReady_3 & (state == 3'h0 | _dpIn_va_T &
    io_in_bits_mixPcMode | _dpIn_va_T_2); // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/Threadgroup.scala 164:41]
  assign io_out_valid = outValid; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/Threadgroup.scala 163:16]
  assign io_out_bits_matrix_d_data = {io_out_bits_matrix_d_data_hi,io_out_bits_matrix_d_data_lo}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/Threadgroup.scala 161:35]
  assign dp_clock = clock;
  assign dp_reset = reset;
  assign dp_io_in_valid = dp_in_valid; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/DotProdUnit.scala 178:20]
  assign dp_io_in_bits_vec_a_0 = _dpIn_va_T_9 | _dpIn_va_T_7; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  assign dp_io_in_bits_vec_a_1 = _dpIn_va_T_16 | _dpIn_va_T_14; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  assign dp_io_in_bits_vec_a_2 = _dpIn_va_T_23 | _dpIn_va_T_21; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  assign dp_io_in_bits_vec_a_3 = _dpIn_va_T_30 | _dpIn_va_T_28; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  assign dp_io_in_bits_vec_b_0 = io_in_bits_matrix_b_data[255:240]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/package.scala 44:28]
  assign dp_io_in_bits_vec_b_1 = io_in_bits_matrix_b_data[239:224]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/package.scala 44:28]
  assign dp_io_in_bits_vec_b_2 = io_in_bits_matrix_b_data[223:208]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/package.scala 44:28]
  assign dp_io_in_bits_vec_b_3 = io_in_bits_matrix_b_data[207:192]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/package.scala 44:28]
  assign dp_io_in_bits_c = _dpIn_c_T_11 | _dpIn_c_T_9; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  assign dp_io_in_bits_mixPc = io_in_bits_mixPcMode; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/DotProdUnit.scala 182:25]
  assign dp_io_in_bits_rowtag = _rowtag_in_T_8 | _rowtag_in_T_6; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  assign dp_1_clock = clock;
  assign dp_1_reset = reset;
  assign dp_1_io_in_valid = dp_in_valid; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/DotProdUnit.scala 178:20]
  assign dp_1_io_in_bits_vec_a_0 = _dpIn_va_T_9 | _dpIn_va_T_7; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  assign dp_1_io_in_bits_vec_a_1 = _dpIn_va_T_16 | _dpIn_va_T_14; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  assign dp_1_io_in_bits_vec_a_2 = _dpIn_va_T_23 | _dpIn_va_T_21; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  assign dp_1_io_in_bits_vec_a_3 = _dpIn_va_T_30 | _dpIn_va_T_28; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  assign dp_1_io_in_bits_vec_b_0 = io_in_bits_matrix_b_data[191:176]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/package.scala 44:28]
  assign dp_1_io_in_bits_vec_b_1 = io_in_bits_matrix_b_data[175:160]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/package.scala 44:28]
  assign dp_1_io_in_bits_vec_b_2 = io_in_bits_matrix_b_data[159:144]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/package.scala 44:28]
  assign dp_1_io_in_bits_vec_b_3 = io_in_bits_matrix_b_data[143:128]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/package.scala 44:28]
  assign dp_1_io_in_bits_c = _dpIn_c_T_18 | _dpIn_c_T_16; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  assign dp_1_io_in_bits_mixPc = io_in_bits_mixPcMode; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/DotProdUnit.scala 182:25]
  assign dp_1_io_in_bits_rowtag = _rowtag_in_T_8 | _rowtag_in_T_6; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  assign dp_2_clock = clock;
  assign dp_2_reset = reset;
  assign dp_2_io_in_valid = dp_in_valid; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/DotProdUnit.scala 178:20]
  assign dp_2_io_in_bits_vec_a_0 = _dpIn_va_T_9 | _dpIn_va_T_7; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  assign dp_2_io_in_bits_vec_a_1 = _dpIn_va_T_16 | _dpIn_va_T_14; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  assign dp_2_io_in_bits_vec_a_2 = _dpIn_va_T_23 | _dpIn_va_T_21; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  assign dp_2_io_in_bits_vec_a_3 = _dpIn_va_T_30 | _dpIn_va_T_28; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  assign dp_2_io_in_bits_vec_b_0 = io_in_bits_matrix_b_data[127:112]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/package.scala 44:28]
  assign dp_2_io_in_bits_vec_b_1 = io_in_bits_matrix_b_data[111:96]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/package.scala 44:28]
  assign dp_2_io_in_bits_vec_b_2 = io_in_bits_matrix_b_data[95:80]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/package.scala 44:28]
  assign dp_2_io_in_bits_vec_b_3 = io_in_bits_matrix_b_data[79:64]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/package.scala 44:28]
  assign dp_2_io_in_bits_c = _dpIn_c_T_25 | _dpIn_c_T_23; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  assign dp_2_io_in_bits_mixPc = io_in_bits_mixPcMode; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/DotProdUnit.scala 182:25]
  assign dp_2_io_in_bits_rowtag = _rowtag_in_T_8 | _rowtag_in_T_6; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  assign dp_3_clock = clock;
  assign dp_3_reset = reset;
  assign dp_3_io_in_valid = dp_in_valid; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/DotProdUnit.scala 178:20]
  assign dp_3_io_in_bits_vec_a_0 = _dpIn_va_T_9 | _dpIn_va_T_7; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  assign dp_3_io_in_bits_vec_a_1 = _dpIn_va_T_16 | _dpIn_va_T_14; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  assign dp_3_io_in_bits_vec_a_2 = _dpIn_va_T_23 | _dpIn_va_T_21; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  assign dp_3_io_in_bits_vec_a_3 = _dpIn_va_T_30 | _dpIn_va_T_28; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  assign dp_3_io_in_bits_vec_b_0 = io_in_bits_matrix_b_data[63:48]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/package.scala 44:28]
  assign dp_3_io_in_bits_vec_b_1 = io_in_bits_matrix_b_data[47:32]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/package.scala 44:28]
  assign dp_3_io_in_bits_vec_b_2 = io_in_bits_matrix_b_data[31:16]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/package.scala 44:28]
  assign dp_3_io_in_bits_vec_b_3 = io_in_bits_matrix_b_data[15:0]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/package.scala 44:28]
  assign dp_3_io_in_bits_c = _dpIn_c_T_32 | _dpIn_c_T_30; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  assign dp_3_io_in_bits_mixPc = io_in_bits_mixPcMode; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/DotProdUnit.scala 182:25]
  assign dp_3_io_in_bits_rowtag = _rowtag_in_T_8 | _rowtag_in_T_6; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  always @(posedge clock) begin
    if (dpValid_0 & dpValid_1 & dpValid_2 & dpValid_3) begin // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/Threadgroup.scala 132:31]
      if (2'h0 == rowtag_out) begin // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/Threadgroup.scala 133:24]
        if (outMixPc) begin // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/Threadgroup.scala 135:24]
          matrix_d_0 <= result_fp32_hi; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/Threadgroup.scala 136:23]
        end else begin
          matrix_d_0 <= result_fp16; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/Threadgroup.scala 139:23]
        end
      end
    end
    if (dpValid_0 & dpValid_1 & dpValid_2 & dpValid_3) begin // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/Threadgroup.scala 132:31]
      if (2'h0 == rowtag_out) begin // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/Threadgroup.scala 133:24]
        if (outMixPc) begin // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/Threadgroup.scala 135:24]
          matrix_d_1 <= result_fp32_lo; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/Threadgroup.scala 137:23]
        end
      end else if (2'h1 == rowtag_out) begin // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/Threadgroup.scala 133:24]
        if (!(outMixPc)) begin // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/Threadgroup.scala 143:24]
          matrix_d_1 <= result_fp16; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/Threadgroup.scala 148:23]
        end
      end
    end
    if (dpValid_0 & dpValid_1 & dpValid_2 & dpValid_3) begin // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/Threadgroup.scala 132:31]
      if (!(2'h0 == rowtag_out)) begin // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/Threadgroup.scala 133:24]
        if (2'h1 == rowtag_out) begin // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/Threadgroup.scala 133:24]
          if (outMixPc) begin // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/Threadgroup.scala 143:24]
            matrix_d_2 <= result_fp32_hi; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/Threadgroup.scala 144:23]
          end
        end else if (2'h2 == rowtag_out) begin // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/Threadgroup.scala 133:24]
          matrix_d_2 <= result_fp16; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/Threadgroup.scala 152:21]
        end
      end
    end
    if (dpValid_0 & dpValid_1 & dpValid_2 & dpValid_3) begin // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/Threadgroup.scala 132:31]
      if (!(2'h0 == rowtag_out)) begin // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/Threadgroup.scala 133:24]
        if (2'h1 == rowtag_out) begin // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/Threadgroup.scala 133:24]
          if (outMixPc) begin // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/Threadgroup.scala 143:24]
            matrix_d_3 <= result_fp32_lo; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/Threadgroup.scala 145:23]
          end
        end else if (!(2'h2 == rowtag_out)) begin // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/Threadgroup.scala 133:24]
          matrix_d_3 <= _GEN_29;
        end
      end
    end
    if (reset) begin // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/Threadgroup.scala 38:25]
      outValid <= 1'h0; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/Threadgroup.scala 38:25]
    end else if (dpValid_0 & dpValid_1 & dpValid_2 & dpValid_3) begin // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/Threadgroup.scala 132:31]
      if (2'h0 == rowtag_out) begin // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/Threadgroup.scala 133:24]
        outValid <= _GEN_0;
      end else if (2'h1 == rowtag_out) begin // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/Threadgroup.scala 133:24]
        outValid <= _GEN_27;
      end else begin
        outValid <= _GEN_33;
      end
    end else begin
      outValid <= _GEN_0;
    end
    if (reset) begin // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/Threadgroup.scala 44:22]
      state <= 3'h0; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/Threadgroup.scala 44:22]
    end else if (3'h0 == state) begin // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/Threadgroup.scala 47:17]
      if (prehandshaked) begin // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/Threadgroup.scala 49:27]
        state <= 3'h1; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/Threadgroup.scala 50:15]
      end
    end else if (3'h1 == state) begin // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/Threadgroup.scala 47:17]
      state <= 3'h2;
    end else if (3'h2 == state) begin // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/Threadgroup.scala 47:17]
      state <= _GEN_6;
    end else begin
      state <= _GEN_15;
    end
    if (reset) begin // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/Threadgroup.scala 45:28]
      dp_in_valid <= 1'h0; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/Threadgroup.scala 45:28]
    end else if (3'h0 == state) begin // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/Threadgroup.scala 47:17]
      dp_in_valid <= prehandshaked;
    end else if (!(3'h1 == state)) begin // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/Threadgroup.scala 47:17]
      if (3'h2 == state) begin // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/Threadgroup.scala 47:17]
        dp_in_valid <= _GEN_7;
      end else begin
        dp_in_valid <= _GEN_16;
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {2{`RANDOM}};
  matrix_d_0 = _RAND_0[63:0];
  _RAND_1 = {2{`RANDOM}};
  matrix_d_1 = _RAND_1[63:0];
  _RAND_2 = {2{`RANDOM}};
  matrix_d_2 = _RAND_2[63:0];
  _RAND_3 = {2{`RANDOM}};
  matrix_d_3 = _RAND_3[63:0];
  _RAND_4 = {1{`RANDOM}};
  outValid = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  state = _RAND_5[2:0];
  _RAND_6 = {1{`RANDOM}};
  dp_in_valid = _RAND_6[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Octet(
  input          clock,
  input          reset,
  output         io_in_ready, // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/Octet.scala 26:14]
  input          io_in_valid, // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/Octet.scala 26:14]
  input  [255:0] io_in_bits_threadgroup0_matrix_a_data, // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/Octet.scala 26:14]
  input  [255:0] io_in_bits_threadgroup0_matrix_b_data, // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/Octet.scala 26:14]
  input  [255:0] io_in_bits_threadgroup0_matrix_c_data, // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/Octet.scala 26:14]
  input  [255:0] io_in_bits_threadgroup4_matrix_a_data, // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/Octet.scala 26:14]
  input  [255:0] io_in_bits_threadgroup4_matrix_b_data, // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/Octet.scala 26:14]
  input  [255:0] io_in_bits_threadgroup4_matrix_c_data, // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/Octet.scala 26:14]
  input          io_in_bits_matBSel, // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/Octet.scala 26:14]
  input          io_in_bits_mixPcMode, // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/Octet.scala 26:14]
  output         io_out_valid, // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/Octet.scala 26:14]
  output [255:0] io_out_bits_threadgroup0_matrix_d_data, // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/Octet.scala 26:14]
  output [255:0] io_out_bits_threadgroup4_matrix_d_data // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/Octet.scala 26:14]
);
  wire  tg_clock; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/Threadgroup.scala 170:20]
  wire  tg_reset; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/Threadgroup.scala 170:20]
  wire  tg_io_in_ready; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/Threadgroup.scala 170:20]
  wire  tg_io_in_valid; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/Threadgroup.scala 170:20]
  wire [255:0] tg_io_in_bits_matrix_a_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/Threadgroup.scala 170:20]
  wire [255:0] tg_io_in_bits_matrix_b_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/Threadgroup.scala 170:20]
  wire [255:0] tg_io_in_bits_matrix_c_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/Threadgroup.scala 170:20]
  wire  tg_io_in_bits_mixPcMode; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/Threadgroup.scala 170:20]
  wire  tg_io_out_valid; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/Threadgroup.scala 170:20]
  wire [255:0] tg_io_out_bits_matrix_d_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/Threadgroup.scala 170:20]
  wire  tg_1_clock; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/Threadgroup.scala 170:20]
  wire  tg_1_reset; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/Threadgroup.scala 170:20]
  wire  tg_1_io_in_ready; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/Threadgroup.scala 170:20]
  wire  tg_1_io_in_valid; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/Threadgroup.scala 170:20]
  wire [255:0] tg_1_io_in_bits_matrix_a_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/Threadgroup.scala 170:20]
  wire [255:0] tg_1_io_in_bits_matrix_b_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/Threadgroup.scala 170:20]
  wire [255:0] tg_1_io_in_bits_matrix_c_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/Threadgroup.scala 170:20]
  wire  tg_1_io_in_bits_mixPcMode; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/Threadgroup.scala 170:20]
  wire  tg_1_io_out_valid; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/Threadgroup.scala 170:20]
  wire [255:0] tg_1_io_out_bits_matrix_d_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/Threadgroup.scala 170:20]
  Threadgroup tg ( // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/Threadgroup.scala 170:20]
    .clock(tg_clock),
    .reset(tg_reset),
    .io_in_ready(tg_io_in_ready),
    .io_in_valid(tg_io_in_valid),
    .io_in_bits_matrix_a_data(tg_io_in_bits_matrix_a_data),
    .io_in_bits_matrix_b_data(tg_io_in_bits_matrix_b_data),
    .io_in_bits_matrix_c_data(tg_io_in_bits_matrix_c_data),
    .io_in_bits_mixPcMode(tg_io_in_bits_mixPcMode),
    .io_out_valid(tg_io_out_valid),
    .io_out_bits_matrix_d_data(tg_io_out_bits_matrix_d_data)
  );
  Threadgroup tg_1 ( // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/Threadgroup.scala 170:20]
    .clock(tg_1_clock),
    .reset(tg_1_reset),
    .io_in_ready(tg_1_io_in_ready),
    .io_in_valid(tg_1_io_in_valid),
    .io_in_bits_matrix_a_data(tg_1_io_in_bits_matrix_a_data),
    .io_in_bits_matrix_b_data(tg_1_io_in_bits_matrix_b_data),
    .io_in_bits_matrix_c_data(tg_1_io_in_bits_matrix_c_data),
    .io_in_bits_mixPcMode(tg_1_io_in_bits_mixPcMode),
    .io_out_valid(tg_1_io_out_valid),
    .io_out_bits_matrix_d_data(tg_1_io_out_bits_matrix_d_data)
  );
  assign io_in_ready = tg_io_in_ready & tg_1_io_in_ready; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/Octet.scala 54:28]
  assign io_out_valid = tg_io_out_valid & tg_1_io_out_valid; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/Octet.scala 55:29]
  assign io_out_bits_threadgroup0_matrix_d_data = tg_io_out_bits_matrix_d_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/Octet.scala 56:37]
  assign io_out_bits_threadgroup4_matrix_d_data = tg_1_io_out_bits_matrix_d_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/Octet.scala 57:37]
  assign tg_clock = clock;
  assign tg_reset = reset;
  assign tg_io_in_valid = io_in_valid; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/Threadgroup.scala 174:20]
  assign tg_io_in_bits_matrix_a_data = io_in_bits_threadgroup0_matrix_a_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/Threadgroup.scala 175:28]
  assign tg_io_in_bits_matrix_b_data = io_in_bits_matBSel ? io_in_bits_threadgroup4_matrix_b_data :
    io_in_bits_threadgroup0_matrix_b_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/Octet.scala 42:22]
  assign tg_io_in_bits_matrix_c_data = io_in_bits_threadgroup0_matrix_c_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/Threadgroup.scala 177:28]
  assign tg_io_in_bits_mixPcMode = io_in_bits_mixPcMode; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/Threadgroup.scala 178:29]
  assign tg_1_clock = clock;
  assign tg_1_reset = reset;
  assign tg_1_io_in_valid = io_in_valid; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/Threadgroup.scala 174:20]
  assign tg_1_io_in_bits_matrix_a_data = io_in_bits_threadgroup4_matrix_a_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/Threadgroup.scala 175:28]
  assign tg_1_io_in_bits_matrix_b_data = io_in_bits_matBSel ? io_in_bits_threadgroup4_matrix_b_data :
    io_in_bits_threadgroup0_matrix_b_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/Octet.scala 45:22]
  assign tg_1_io_in_bits_matrix_c_data = io_in_bits_threadgroup4_matrix_c_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/Threadgroup.scala 177:28]
  assign tg_1_io_in_bits_mixPcMode = io_in_bits_mixPcMode; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/Threadgroup.scala 178:29]
endmodule
module TensorCore(
  input          clock,
  input          reset,
  output         io_in_ready, // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/TensorCore.scala 26:14]
  input          io_in_valid, // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/TensorCore.scala 26:14]
  input  [255:0] io_in_bits_octet0_threadgroup0_matrix_a_data, // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/TensorCore.scala 26:14]
  input  [255:0] io_in_bits_octet0_threadgroup0_matrix_b_data, // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/TensorCore.scala 26:14]
  input  [255:0] io_in_bits_octet0_threadgroup0_matrix_c_data, // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/TensorCore.scala 26:14]
  input  [255:0] io_in_bits_octet0_threadgroup4_matrix_a_data, // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/TensorCore.scala 26:14]
  input  [255:0] io_in_bits_octet0_threadgroup4_matrix_b_data, // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/TensorCore.scala 26:14]
  input  [255:0] io_in_bits_octet0_threadgroup4_matrix_c_data, // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/TensorCore.scala 26:14]
  input  [255:0] io_in_bits_octet1_threadgroup0_matrix_a_data, // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/TensorCore.scala 26:14]
  input  [255:0] io_in_bits_octet1_threadgroup0_matrix_b_data, // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/TensorCore.scala 26:14]
  input  [255:0] io_in_bits_octet1_threadgroup0_matrix_c_data, // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/TensorCore.scala 26:14]
  input  [255:0] io_in_bits_octet1_threadgroup4_matrix_a_data, // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/TensorCore.scala 26:14]
  input  [255:0] io_in_bits_octet1_threadgroup4_matrix_b_data, // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/TensorCore.scala 26:14]
  input  [255:0] io_in_bits_octet1_threadgroup4_matrix_c_data, // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/TensorCore.scala 26:14]
  input          io_in_bits_ctrl_matBSel, // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/TensorCore.scala 26:14]
  input          io_in_bits_ctrl_mixPcMode, // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/TensorCore.scala 26:14]
  output         io_out_valid, // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/TensorCore.scala 26:14]
  output [255:0] io_out_bits_octet0_threadgroup0_matrix_d_data, // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/TensorCore.scala 26:14]
  output [255:0] io_out_bits_octet0_threadgroup4_matrix_d_data, // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/TensorCore.scala 26:14]
  output [255:0] io_out_bits_octet1_threadgroup0_matrix_d_data, // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/TensorCore.scala 26:14]
  output [255:0] io_out_bits_octet1_threadgroup4_matrix_d_data // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/TensorCore.scala 26:14]
);
  wire  ot_clock; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/Octet.scala 66:20]
  wire  ot_reset; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/Octet.scala 66:20]
  wire  ot_io_in_ready; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/Octet.scala 66:20]
  wire  ot_io_in_valid; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/Octet.scala 66:20]
  wire [255:0] ot_io_in_bits_threadgroup0_matrix_a_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/Octet.scala 66:20]
  wire [255:0] ot_io_in_bits_threadgroup0_matrix_b_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/Octet.scala 66:20]
  wire [255:0] ot_io_in_bits_threadgroup0_matrix_c_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/Octet.scala 66:20]
  wire [255:0] ot_io_in_bits_threadgroup4_matrix_a_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/Octet.scala 66:20]
  wire [255:0] ot_io_in_bits_threadgroup4_matrix_b_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/Octet.scala 66:20]
  wire [255:0] ot_io_in_bits_threadgroup4_matrix_c_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/Octet.scala 66:20]
  wire  ot_io_in_bits_matBSel; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/Octet.scala 66:20]
  wire  ot_io_in_bits_mixPcMode; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/Octet.scala 66:20]
  wire  ot_io_out_valid; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/Octet.scala 66:20]
  wire [255:0] ot_io_out_bits_threadgroup0_matrix_d_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/Octet.scala 66:20]
  wire [255:0] ot_io_out_bits_threadgroup4_matrix_d_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/Octet.scala 66:20]
  wire  ot_1_clock; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/Octet.scala 66:20]
  wire  ot_1_reset; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/Octet.scala 66:20]
  wire  ot_1_io_in_ready; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/Octet.scala 66:20]
  wire  ot_1_io_in_valid; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/Octet.scala 66:20]
  wire [255:0] ot_1_io_in_bits_threadgroup0_matrix_a_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/Octet.scala 66:20]
  wire [255:0] ot_1_io_in_bits_threadgroup0_matrix_b_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/Octet.scala 66:20]
  wire [255:0] ot_1_io_in_bits_threadgroup0_matrix_c_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/Octet.scala 66:20]
  wire [255:0] ot_1_io_in_bits_threadgroup4_matrix_a_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/Octet.scala 66:20]
  wire [255:0] ot_1_io_in_bits_threadgroup4_matrix_b_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/Octet.scala 66:20]
  wire [255:0] ot_1_io_in_bits_threadgroup4_matrix_c_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/Octet.scala 66:20]
  wire  ot_1_io_in_bits_matBSel; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/Octet.scala 66:20]
  wire  ot_1_io_in_bits_mixPcMode; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/Octet.scala 66:20]
  wire  ot_1_io_out_valid; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/Octet.scala 66:20]
  wire [255:0] ot_1_io_out_bits_threadgroup0_matrix_d_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/Octet.scala 66:20]
  wire [255:0] ot_1_io_out_bits_threadgroup4_matrix_d_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/Octet.scala 66:20]
  wire  ot_ready_0 = ot_io_in_ready; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/TensorCore.scala 41:22 48:17]
  wire  ot_ready_1 = ot_1_io_in_ready; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/TensorCore.scala 41:22 48:17]
  wire  ot_valid_0 = ot_io_out_valid; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/TensorCore.scala 40:22 47:17]
  wire  ot_valid_1 = ot_1_io_out_valid; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/TensorCore.scala 40:22 47:17]
  Octet ot ( // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/Octet.scala 66:20]
    .clock(ot_clock),
    .reset(ot_reset),
    .io_in_ready(ot_io_in_ready),
    .io_in_valid(ot_io_in_valid),
    .io_in_bits_threadgroup0_matrix_a_data(ot_io_in_bits_threadgroup0_matrix_a_data),
    .io_in_bits_threadgroup0_matrix_b_data(ot_io_in_bits_threadgroup0_matrix_b_data),
    .io_in_bits_threadgroup0_matrix_c_data(ot_io_in_bits_threadgroup0_matrix_c_data),
    .io_in_bits_threadgroup4_matrix_a_data(ot_io_in_bits_threadgroup4_matrix_a_data),
    .io_in_bits_threadgroup4_matrix_b_data(ot_io_in_bits_threadgroup4_matrix_b_data),
    .io_in_bits_threadgroup4_matrix_c_data(ot_io_in_bits_threadgroup4_matrix_c_data),
    .io_in_bits_matBSel(ot_io_in_bits_matBSel),
    .io_in_bits_mixPcMode(ot_io_in_bits_mixPcMode),
    .io_out_valid(ot_io_out_valid),
    .io_out_bits_threadgroup0_matrix_d_data(ot_io_out_bits_threadgroup0_matrix_d_data),
    .io_out_bits_threadgroup4_matrix_d_data(ot_io_out_bits_threadgroup4_matrix_d_data)
  );
  Octet ot_1 ( // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/Octet.scala 66:20]
    .clock(ot_1_clock),
    .reset(ot_1_reset),
    .io_in_ready(ot_1_io_in_ready),
    .io_in_valid(ot_1_io_in_valid),
    .io_in_bits_threadgroup0_matrix_a_data(ot_1_io_in_bits_threadgroup0_matrix_a_data),
    .io_in_bits_threadgroup0_matrix_b_data(ot_1_io_in_bits_threadgroup0_matrix_b_data),
    .io_in_bits_threadgroup0_matrix_c_data(ot_1_io_in_bits_threadgroup0_matrix_c_data),
    .io_in_bits_threadgroup4_matrix_a_data(ot_1_io_in_bits_threadgroup4_matrix_a_data),
    .io_in_bits_threadgroup4_matrix_b_data(ot_1_io_in_bits_threadgroup4_matrix_b_data),
    .io_in_bits_threadgroup4_matrix_c_data(ot_1_io_in_bits_threadgroup4_matrix_c_data),
    .io_in_bits_matBSel(ot_1_io_in_bits_matBSel),
    .io_in_bits_mixPcMode(ot_1_io_in_bits_mixPcMode),
    .io_out_valid(ot_1_io_out_valid),
    .io_out_bits_threadgroup0_matrix_d_data(ot_1_io_out_bits_threadgroup0_matrix_d_data),
    .io_out_bits_threadgroup4_matrix_d_data(ot_1_io_out_bits_threadgroup4_matrix_d_data)
  );
  assign io_in_ready = ot_ready_0 & ot_ready_1; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/TensorCore.scala 51:36]
  assign io_out_valid = ot_valid_0 & ot_valid_1; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/TensorCore.scala 52:36]
  assign io_out_bits_octet0_threadgroup0_matrix_d_data = ot_io_out_bits_threadgroup0_matrix_d_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/TensorCore.scala 46:{27,27}]
  assign io_out_bits_octet0_threadgroup4_matrix_d_data = ot_io_out_bits_threadgroup4_matrix_d_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/TensorCore.scala 46:{27,27}]
  assign io_out_bits_octet1_threadgroup0_matrix_d_data = ot_1_io_out_bits_threadgroup0_matrix_d_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/TensorCore.scala 46:{27,27}]
  assign io_out_bits_octet1_threadgroup4_matrix_d_data = ot_1_io_out_bits_threadgroup4_matrix_d_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/TensorCore.scala 46:{27,27}]
  assign ot_clock = clock;
  assign ot_reset = reset;
  assign ot_io_in_valid = io_in_valid; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/Octet.scala 77:20]
  assign ot_io_in_bits_threadgroup0_matrix_a_data = io_in_bits_octet0_threadgroup0_matrix_a_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/TensorCore.scala 37:{22,22}]
  assign ot_io_in_bits_threadgroup0_matrix_b_data = io_in_bits_octet0_threadgroup0_matrix_b_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/TensorCore.scala 37:{22,22}]
  assign ot_io_in_bits_threadgroup0_matrix_c_data = io_in_bits_octet0_threadgroup0_matrix_c_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/TensorCore.scala 37:{22,22}]
  assign ot_io_in_bits_threadgroup4_matrix_a_data = io_in_bits_octet0_threadgroup4_matrix_a_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/TensorCore.scala 37:{22,22}]
  assign ot_io_in_bits_threadgroup4_matrix_b_data = io_in_bits_octet0_threadgroup4_matrix_b_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/TensorCore.scala 37:{22,22}]
  assign ot_io_in_bits_threadgroup4_matrix_c_data = io_in_bits_octet0_threadgroup4_matrix_c_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/TensorCore.scala 37:{22,22}]
  assign ot_io_in_bits_matBSel = io_in_bits_ctrl_matBSel; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/Octet.scala 84:27]
  assign ot_io_in_bits_mixPcMode = io_in_bits_ctrl_mixPcMode; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/Octet.scala 85:29]
  assign ot_1_clock = clock;
  assign ot_1_reset = reset;
  assign ot_1_io_in_valid = io_in_valid; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/Octet.scala 77:20]
  assign ot_1_io_in_bits_threadgroup0_matrix_a_data = io_in_bits_octet1_threadgroup0_matrix_a_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/TensorCore.scala 37:{22,22}]
  assign ot_1_io_in_bits_threadgroup0_matrix_b_data = io_in_bits_octet1_threadgroup0_matrix_b_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/TensorCore.scala 37:{22,22}]
  assign ot_1_io_in_bits_threadgroup0_matrix_c_data = io_in_bits_octet1_threadgroup0_matrix_c_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/TensorCore.scala 37:{22,22}]
  assign ot_1_io_in_bits_threadgroup4_matrix_a_data = io_in_bits_octet1_threadgroup4_matrix_a_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/TensorCore.scala 37:{22,22}]
  assign ot_1_io_in_bits_threadgroup4_matrix_b_data = io_in_bits_octet1_threadgroup4_matrix_b_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/TensorCore.scala 37:{22,22}]
  assign ot_1_io_in_bits_threadgroup4_matrix_c_data = io_in_bits_octet1_threadgroup4_matrix_c_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/TensorCore.scala 37:{22,22}]
  assign ot_1_io_in_bits_matBSel = io_in_bits_ctrl_matBSel; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/Octet.scala 84:27]
  assign ot_1_io_in_bits_mixPcMode = io_in_bits_ctrl_mixPcMode; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/Octet.scala 85:29]
endmodule
module Top(
  input          clock,
  input          reset,
  output         io_in_ready, // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/Top.scala 43:14]
  input          io_in_valid, // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/Top.scala 43:14]
  input  [255:0] io_in_bits_tc0_ot0_tg0_matrix_a, // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/Top.scala 43:14]
  input  [255:0] io_in_bits_tc0_ot0_tg0_matrix_b, // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/Top.scala 43:14]
  input  [255:0] io_in_bits_tc0_ot0_tg0_matrix_c, // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/Top.scala 43:14]
  input  [255:0] io_in_bits_tc0_ot0_tg4_matrix_a, // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/Top.scala 43:14]
  input  [255:0] io_in_bits_tc0_ot0_tg4_matrix_b, // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/Top.scala 43:14]
  input  [255:0] io_in_bits_tc0_ot0_tg4_matrix_c, // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/Top.scala 43:14]
  input  [255:0] io_in_bits_tc0_ot1_tg0_matrix_a, // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/Top.scala 43:14]
  input  [255:0] io_in_bits_tc0_ot1_tg0_matrix_b, // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/Top.scala 43:14]
  input  [255:0] io_in_bits_tc0_ot1_tg0_matrix_c, // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/Top.scala 43:14]
  input  [255:0] io_in_bits_tc0_ot1_tg4_matrix_a, // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/Top.scala 43:14]
  input  [255:0] io_in_bits_tc0_ot1_tg4_matrix_b, // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/Top.scala 43:14]
  input  [255:0] io_in_bits_tc0_ot1_tg4_matrix_c, // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/Top.scala 43:14]
  input  [255:0] io_in_bits_tc1_ot0_tg0_matrix_a, // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/Top.scala 43:14]
  input  [255:0] io_in_bits_tc1_ot0_tg0_matrix_b, // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/Top.scala 43:14]
  input  [255:0] io_in_bits_tc1_ot0_tg0_matrix_c, // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/Top.scala 43:14]
  input  [255:0] io_in_bits_tc1_ot0_tg4_matrix_a, // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/Top.scala 43:14]
  input  [255:0] io_in_bits_tc1_ot0_tg4_matrix_b, // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/Top.scala 43:14]
  input  [255:0] io_in_bits_tc1_ot0_tg4_matrix_c, // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/Top.scala 43:14]
  input  [255:0] io_in_bits_tc1_ot1_tg0_matrix_a, // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/Top.scala 43:14]
  input  [255:0] io_in_bits_tc1_ot1_tg0_matrix_b, // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/Top.scala 43:14]
  input  [255:0] io_in_bits_tc1_ot1_tg0_matrix_c, // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/Top.scala 43:14]
  input  [255:0] io_in_bits_tc1_ot1_tg4_matrix_a, // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/Top.scala 43:14]
  input  [255:0] io_in_bits_tc1_ot1_tg4_matrix_b, // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/Top.scala 43:14]
  input  [255:0] io_in_bits_tc1_ot1_tg4_matrix_c, // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/Top.scala 43:14]
  input          io_in_bits_ctrl_matBSel, // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/Top.scala 43:14]
  input          io_in_bits_ctrl_mixPcMode, // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/Top.scala 43:14]
  output         io_out_valid, // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/Top.scala 43:14]
  output [255:0] io_out_bits_tc0_octet0_threadgroup0_matrix_d_data, // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/Top.scala 43:14]
  output [255:0] io_out_bits_tc0_octet0_threadgroup4_matrix_d_data, // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/Top.scala 43:14]
  output [255:0] io_out_bits_tc0_octet1_threadgroup0_matrix_d_data, // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/Top.scala 43:14]
  output [255:0] io_out_bits_tc0_octet1_threadgroup4_matrix_d_data, // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/Top.scala 43:14]
  output [255:0] io_out_bits_tc1_octet0_threadgroup0_matrix_d_data, // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/Top.scala 43:14]
  output [255:0] io_out_bits_tc1_octet0_threadgroup4_matrix_d_data, // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/Top.scala 43:14]
  output [255:0] io_out_bits_tc1_octet1_threadgroup0_matrix_d_data, // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/Top.scala 43:14]
  output [255:0] io_out_bits_tc1_octet1_threadgroup4_matrix_d_data // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/Top.scala 43:14]
);
  wire  tc_clock; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/TensorCore.scala 67:20]
  wire  tc_reset; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/TensorCore.scala 67:20]
  wire  tc_io_in_ready; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/TensorCore.scala 67:20]
  wire  tc_io_in_valid; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/TensorCore.scala 67:20]
  wire [255:0] tc_io_in_bits_octet0_threadgroup0_matrix_a_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/TensorCore.scala 67:20]
  wire [255:0] tc_io_in_bits_octet0_threadgroup0_matrix_b_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/TensorCore.scala 67:20]
  wire [255:0] tc_io_in_bits_octet0_threadgroup0_matrix_c_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/TensorCore.scala 67:20]
  wire [255:0] tc_io_in_bits_octet0_threadgroup4_matrix_a_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/TensorCore.scala 67:20]
  wire [255:0] tc_io_in_bits_octet0_threadgroup4_matrix_b_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/TensorCore.scala 67:20]
  wire [255:0] tc_io_in_bits_octet0_threadgroup4_matrix_c_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/TensorCore.scala 67:20]
  wire [255:0] tc_io_in_bits_octet1_threadgroup0_matrix_a_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/TensorCore.scala 67:20]
  wire [255:0] tc_io_in_bits_octet1_threadgroup0_matrix_b_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/TensorCore.scala 67:20]
  wire [255:0] tc_io_in_bits_octet1_threadgroup0_matrix_c_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/TensorCore.scala 67:20]
  wire [255:0] tc_io_in_bits_octet1_threadgroup4_matrix_a_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/TensorCore.scala 67:20]
  wire [255:0] tc_io_in_bits_octet1_threadgroup4_matrix_b_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/TensorCore.scala 67:20]
  wire [255:0] tc_io_in_bits_octet1_threadgroup4_matrix_c_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/TensorCore.scala 67:20]
  wire  tc_io_in_bits_ctrl_matBSel; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/TensorCore.scala 67:20]
  wire  tc_io_in_bits_ctrl_mixPcMode; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/TensorCore.scala 67:20]
  wire  tc_io_out_valid; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/TensorCore.scala 67:20]
  wire [255:0] tc_io_out_bits_octet0_threadgroup0_matrix_d_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/TensorCore.scala 67:20]
  wire [255:0] tc_io_out_bits_octet0_threadgroup4_matrix_d_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/TensorCore.scala 67:20]
  wire [255:0] tc_io_out_bits_octet1_threadgroup0_matrix_d_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/TensorCore.scala 67:20]
  wire [255:0] tc_io_out_bits_octet1_threadgroup4_matrix_d_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/TensorCore.scala 67:20]
  wire  tc_1_clock; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/TensorCore.scala 67:20]
  wire  tc_1_reset; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/TensorCore.scala 67:20]
  wire  tc_1_io_in_ready; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/TensorCore.scala 67:20]
  wire  tc_1_io_in_valid; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/TensorCore.scala 67:20]
  wire [255:0] tc_1_io_in_bits_octet0_threadgroup0_matrix_a_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/TensorCore.scala 67:20]
  wire [255:0] tc_1_io_in_bits_octet0_threadgroup0_matrix_b_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/TensorCore.scala 67:20]
  wire [255:0] tc_1_io_in_bits_octet0_threadgroup0_matrix_c_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/TensorCore.scala 67:20]
  wire [255:0] tc_1_io_in_bits_octet0_threadgroup4_matrix_a_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/TensorCore.scala 67:20]
  wire [255:0] tc_1_io_in_bits_octet0_threadgroup4_matrix_b_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/TensorCore.scala 67:20]
  wire [255:0] tc_1_io_in_bits_octet0_threadgroup4_matrix_c_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/TensorCore.scala 67:20]
  wire [255:0] tc_1_io_in_bits_octet1_threadgroup0_matrix_a_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/TensorCore.scala 67:20]
  wire [255:0] tc_1_io_in_bits_octet1_threadgroup0_matrix_b_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/TensorCore.scala 67:20]
  wire [255:0] tc_1_io_in_bits_octet1_threadgroup0_matrix_c_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/TensorCore.scala 67:20]
  wire [255:0] tc_1_io_in_bits_octet1_threadgroup4_matrix_a_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/TensorCore.scala 67:20]
  wire [255:0] tc_1_io_in_bits_octet1_threadgroup4_matrix_b_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/TensorCore.scala 67:20]
  wire [255:0] tc_1_io_in_bits_octet1_threadgroup4_matrix_c_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/TensorCore.scala 67:20]
  wire  tc_1_io_in_bits_ctrl_matBSel; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/TensorCore.scala 67:20]
  wire  tc_1_io_in_bits_ctrl_mixPcMode; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/TensorCore.scala 67:20]
  wire  tc_1_io_out_valid; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/TensorCore.scala 67:20]
  wire [255:0] tc_1_io_out_bits_octet0_threadgroup0_matrix_d_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/TensorCore.scala 67:20]
  wire [255:0] tc_1_io_out_bits_octet0_threadgroup4_matrix_d_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/TensorCore.scala 67:20]
  wire [255:0] tc_1_io_out_bits_octet1_threadgroup0_matrix_d_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/TensorCore.scala 67:20]
  wire [255:0] tc_1_io_out_bits_octet1_threadgroup4_matrix_d_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/TensorCore.scala 67:20]
  wire [15:0] ot0_tg0_matrix_b_matVType__0_0 = io_in_bits_tc0_ot0_tg0_matrix_b[255:240]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/package.scala 77:32]
  wire [15:0] ot0_tg0_matrix_b_matVType__0_1 = io_in_bits_tc0_ot0_tg0_matrix_b[239:224]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/package.scala 77:32]
  wire [15:0] ot0_tg0_matrix_b_matVType__0_2 = io_in_bits_tc0_ot0_tg0_matrix_b[223:208]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/package.scala 77:32]
  wire [15:0] ot0_tg0_matrix_b_matVType__0_3 = io_in_bits_tc0_ot0_tg0_matrix_b[207:192]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/package.scala 77:32]
  wire [15:0] ot0_tg0_matrix_b_matVType__1_0 = io_in_bits_tc0_ot0_tg0_matrix_b[191:176]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/package.scala 77:32]
  wire [15:0] ot0_tg0_matrix_b_matVType__1_1 = io_in_bits_tc0_ot0_tg0_matrix_b[175:160]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/package.scala 77:32]
  wire [15:0] ot0_tg0_matrix_b_matVType__1_2 = io_in_bits_tc0_ot0_tg0_matrix_b[159:144]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/package.scala 77:32]
  wire [15:0] ot0_tg0_matrix_b_matVType__1_3 = io_in_bits_tc0_ot0_tg0_matrix_b[143:128]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/package.scala 77:32]
  wire [15:0] ot0_tg0_matrix_b_matVType__2_0 = io_in_bits_tc0_ot0_tg0_matrix_b[127:112]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/package.scala 77:32]
  wire [15:0] ot0_tg0_matrix_b_matVType__2_1 = io_in_bits_tc0_ot0_tg0_matrix_b[111:96]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/package.scala 77:32]
  wire [15:0] ot0_tg0_matrix_b_matVType__2_2 = io_in_bits_tc0_ot0_tg0_matrix_b[95:80]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/package.scala 77:32]
  wire [15:0] ot0_tg0_matrix_b_matVType__2_3 = io_in_bits_tc0_ot0_tg0_matrix_b[79:64]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/package.scala 77:32]
  wire [15:0] ot0_tg0_matrix_b_matVType__3_0 = io_in_bits_tc0_ot0_tg0_matrix_b[63:48]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/package.scala 77:32]
  wire [15:0] ot0_tg0_matrix_b_matVType__3_1 = io_in_bits_tc0_ot0_tg0_matrix_b[47:32]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/package.scala 77:32]
  wire [15:0] ot0_tg0_matrix_b_matVType__3_2 = io_in_bits_tc0_ot0_tg0_matrix_b[31:16]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/package.scala 77:32]
  wire [15:0] ot0_tg0_matrix_b_matVType__3_3 = io_in_bits_tc0_ot0_tg0_matrix_b[15:0]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/package.scala 77:32]
  wire [127:0] ot0_tg0_matrix_b_mat_data_lo = {ot0_tg0_matrix_b_matVType__0_2,ot0_tg0_matrix_b_matVType__1_2,
    ot0_tg0_matrix_b_matVType__2_2,ot0_tg0_matrix_b_matVType__3_2,ot0_tg0_matrix_b_matVType__0_3,
    ot0_tg0_matrix_b_matVType__1_3,ot0_tg0_matrix_b_matVType__2_3,ot0_tg0_matrix_b_matVType__3_3}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/package.scala 80:41]
  wire [127:0] ot0_tg0_matrix_b_mat_data_hi = {ot0_tg0_matrix_b_matVType__0_0,ot0_tg0_matrix_b_matVType__1_0,
    ot0_tg0_matrix_b_matVType__2_0,ot0_tg0_matrix_b_matVType__3_0,ot0_tg0_matrix_b_matVType__0_1,
    ot0_tg0_matrix_b_matVType__1_1,ot0_tg0_matrix_b_matVType__2_1,ot0_tg0_matrix_b_matVType__3_1}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/package.scala 80:41]
  wire [15:0] ot0_tg4_matrix_b_matVType__0_0 = io_in_bits_tc0_ot0_tg4_matrix_b[255:240]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/package.scala 77:32]
  wire [15:0] ot0_tg4_matrix_b_matVType__0_1 = io_in_bits_tc0_ot0_tg4_matrix_b[239:224]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/package.scala 77:32]
  wire [15:0] ot0_tg4_matrix_b_matVType__0_2 = io_in_bits_tc0_ot0_tg4_matrix_b[223:208]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/package.scala 77:32]
  wire [15:0] ot0_tg4_matrix_b_matVType__0_3 = io_in_bits_tc0_ot0_tg4_matrix_b[207:192]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/package.scala 77:32]
  wire [15:0] ot0_tg4_matrix_b_matVType__1_0 = io_in_bits_tc0_ot0_tg4_matrix_b[191:176]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/package.scala 77:32]
  wire [15:0] ot0_tg4_matrix_b_matVType__1_1 = io_in_bits_tc0_ot0_tg4_matrix_b[175:160]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/package.scala 77:32]
  wire [15:0] ot0_tg4_matrix_b_matVType__1_2 = io_in_bits_tc0_ot0_tg4_matrix_b[159:144]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/package.scala 77:32]
  wire [15:0] ot0_tg4_matrix_b_matVType__1_3 = io_in_bits_tc0_ot0_tg4_matrix_b[143:128]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/package.scala 77:32]
  wire [15:0] ot0_tg4_matrix_b_matVType__2_0 = io_in_bits_tc0_ot0_tg4_matrix_b[127:112]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/package.scala 77:32]
  wire [15:0] ot0_tg4_matrix_b_matVType__2_1 = io_in_bits_tc0_ot0_tg4_matrix_b[111:96]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/package.scala 77:32]
  wire [15:0] ot0_tg4_matrix_b_matVType__2_2 = io_in_bits_tc0_ot0_tg4_matrix_b[95:80]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/package.scala 77:32]
  wire [15:0] ot0_tg4_matrix_b_matVType__2_3 = io_in_bits_tc0_ot0_tg4_matrix_b[79:64]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/package.scala 77:32]
  wire [15:0] ot0_tg4_matrix_b_matVType__3_0 = io_in_bits_tc0_ot0_tg4_matrix_b[63:48]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/package.scala 77:32]
  wire [15:0] ot0_tg4_matrix_b_matVType__3_1 = io_in_bits_tc0_ot0_tg4_matrix_b[47:32]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/package.scala 77:32]
  wire [15:0] ot0_tg4_matrix_b_matVType__3_2 = io_in_bits_tc0_ot0_tg4_matrix_b[31:16]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/package.scala 77:32]
  wire [15:0] ot0_tg4_matrix_b_matVType__3_3 = io_in_bits_tc0_ot0_tg4_matrix_b[15:0]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/package.scala 77:32]
  wire [127:0] ot0_tg4_matrix_b_mat_data_lo = {ot0_tg4_matrix_b_matVType__0_2,ot0_tg4_matrix_b_matVType__1_2,
    ot0_tg4_matrix_b_matVType__2_2,ot0_tg4_matrix_b_matVType__3_2,ot0_tg4_matrix_b_matVType__0_3,
    ot0_tg4_matrix_b_matVType__1_3,ot0_tg4_matrix_b_matVType__2_3,ot0_tg4_matrix_b_matVType__3_3}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/package.scala 80:41]
  wire [127:0] ot0_tg4_matrix_b_mat_data_hi = {ot0_tg4_matrix_b_matVType__0_0,ot0_tg4_matrix_b_matVType__1_0,
    ot0_tg4_matrix_b_matVType__2_0,ot0_tg4_matrix_b_matVType__3_0,ot0_tg4_matrix_b_matVType__0_1,
    ot0_tg4_matrix_b_matVType__1_1,ot0_tg4_matrix_b_matVType__2_1,ot0_tg4_matrix_b_matVType__3_1}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/package.scala 80:41]
  wire [15:0] ot1_tg0_matrix_b_matVType__0_0 = io_in_bits_tc0_ot1_tg0_matrix_b[255:240]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/package.scala 77:32]
  wire [15:0] ot1_tg0_matrix_b_matVType__0_1 = io_in_bits_tc0_ot1_tg0_matrix_b[239:224]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/package.scala 77:32]
  wire [15:0] ot1_tg0_matrix_b_matVType__0_2 = io_in_bits_tc0_ot1_tg0_matrix_b[223:208]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/package.scala 77:32]
  wire [15:0] ot1_tg0_matrix_b_matVType__0_3 = io_in_bits_tc0_ot1_tg0_matrix_b[207:192]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/package.scala 77:32]
  wire [15:0] ot1_tg0_matrix_b_matVType__1_0 = io_in_bits_tc0_ot1_tg0_matrix_b[191:176]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/package.scala 77:32]
  wire [15:0] ot1_tg0_matrix_b_matVType__1_1 = io_in_bits_tc0_ot1_tg0_matrix_b[175:160]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/package.scala 77:32]
  wire [15:0] ot1_tg0_matrix_b_matVType__1_2 = io_in_bits_tc0_ot1_tg0_matrix_b[159:144]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/package.scala 77:32]
  wire [15:0] ot1_tg0_matrix_b_matVType__1_3 = io_in_bits_tc0_ot1_tg0_matrix_b[143:128]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/package.scala 77:32]
  wire [15:0] ot1_tg0_matrix_b_matVType__2_0 = io_in_bits_tc0_ot1_tg0_matrix_b[127:112]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/package.scala 77:32]
  wire [15:0] ot1_tg0_matrix_b_matVType__2_1 = io_in_bits_tc0_ot1_tg0_matrix_b[111:96]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/package.scala 77:32]
  wire [15:0] ot1_tg0_matrix_b_matVType__2_2 = io_in_bits_tc0_ot1_tg0_matrix_b[95:80]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/package.scala 77:32]
  wire [15:0] ot1_tg0_matrix_b_matVType__2_3 = io_in_bits_tc0_ot1_tg0_matrix_b[79:64]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/package.scala 77:32]
  wire [15:0] ot1_tg0_matrix_b_matVType__3_0 = io_in_bits_tc0_ot1_tg0_matrix_b[63:48]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/package.scala 77:32]
  wire [15:0] ot1_tg0_matrix_b_matVType__3_1 = io_in_bits_tc0_ot1_tg0_matrix_b[47:32]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/package.scala 77:32]
  wire [15:0] ot1_tg0_matrix_b_matVType__3_2 = io_in_bits_tc0_ot1_tg0_matrix_b[31:16]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/package.scala 77:32]
  wire [15:0] ot1_tg0_matrix_b_matVType__3_3 = io_in_bits_tc0_ot1_tg0_matrix_b[15:0]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/package.scala 77:32]
  wire [127:0] ot1_tg0_matrix_b_mat_data_lo = {ot1_tg0_matrix_b_matVType__0_2,ot1_tg0_matrix_b_matVType__1_2,
    ot1_tg0_matrix_b_matVType__2_2,ot1_tg0_matrix_b_matVType__3_2,ot1_tg0_matrix_b_matVType__0_3,
    ot1_tg0_matrix_b_matVType__1_3,ot1_tg0_matrix_b_matVType__2_3,ot1_tg0_matrix_b_matVType__3_3}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/package.scala 80:41]
  wire [127:0] ot1_tg0_matrix_b_mat_data_hi = {ot1_tg0_matrix_b_matVType__0_0,ot1_tg0_matrix_b_matVType__1_0,
    ot1_tg0_matrix_b_matVType__2_0,ot1_tg0_matrix_b_matVType__3_0,ot1_tg0_matrix_b_matVType__0_1,
    ot1_tg0_matrix_b_matVType__1_1,ot1_tg0_matrix_b_matVType__2_1,ot1_tg0_matrix_b_matVType__3_1}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/package.scala 80:41]
  wire [15:0] ot1_tg4_matrix_b_matVType__0_0 = io_in_bits_tc0_ot1_tg4_matrix_b[255:240]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/package.scala 77:32]
  wire [15:0] ot1_tg4_matrix_b_matVType__0_1 = io_in_bits_tc0_ot1_tg4_matrix_b[239:224]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/package.scala 77:32]
  wire [15:0] ot1_tg4_matrix_b_matVType__0_2 = io_in_bits_tc0_ot1_tg4_matrix_b[223:208]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/package.scala 77:32]
  wire [15:0] ot1_tg4_matrix_b_matVType__0_3 = io_in_bits_tc0_ot1_tg4_matrix_b[207:192]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/package.scala 77:32]
  wire [15:0] ot1_tg4_matrix_b_matVType__1_0 = io_in_bits_tc0_ot1_tg4_matrix_b[191:176]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/package.scala 77:32]
  wire [15:0] ot1_tg4_matrix_b_matVType__1_1 = io_in_bits_tc0_ot1_tg4_matrix_b[175:160]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/package.scala 77:32]
  wire [15:0] ot1_tg4_matrix_b_matVType__1_2 = io_in_bits_tc0_ot1_tg4_matrix_b[159:144]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/package.scala 77:32]
  wire [15:0] ot1_tg4_matrix_b_matVType__1_3 = io_in_bits_tc0_ot1_tg4_matrix_b[143:128]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/package.scala 77:32]
  wire [15:0] ot1_tg4_matrix_b_matVType__2_0 = io_in_bits_tc0_ot1_tg4_matrix_b[127:112]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/package.scala 77:32]
  wire [15:0] ot1_tg4_matrix_b_matVType__2_1 = io_in_bits_tc0_ot1_tg4_matrix_b[111:96]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/package.scala 77:32]
  wire [15:0] ot1_tg4_matrix_b_matVType__2_2 = io_in_bits_tc0_ot1_tg4_matrix_b[95:80]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/package.scala 77:32]
  wire [15:0] ot1_tg4_matrix_b_matVType__2_3 = io_in_bits_tc0_ot1_tg4_matrix_b[79:64]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/package.scala 77:32]
  wire [15:0] ot1_tg4_matrix_b_matVType__3_0 = io_in_bits_tc0_ot1_tg4_matrix_b[63:48]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/package.scala 77:32]
  wire [15:0] ot1_tg4_matrix_b_matVType__3_1 = io_in_bits_tc0_ot1_tg4_matrix_b[47:32]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/package.scala 77:32]
  wire [15:0] ot1_tg4_matrix_b_matVType__3_2 = io_in_bits_tc0_ot1_tg4_matrix_b[31:16]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/package.scala 77:32]
  wire [15:0] ot1_tg4_matrix_b_matVType__3_3 = io_in_bits_tc0_ot1_tg4_matrix_b[15:0]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/package.scala 77:32]
  wire [127:0] ot1_tg4_matrix_b_mat_data_lo = {ot1_tg4_matrix_b_matVType__0_2,ot1_tg4_matrix_b_matVType__1_2,
    ot1_tg4_matrix_b_matVType__2_2,ot1_tg4_matrix_b_matVType__3_2,ot1_tg4_matrix_b_matVType__0_3,
    ot1_tg4_matrix_b_matVType__1_3,ot1_tg4_matrix_b_matVType__2_3,ot1_tg4_matrix_b_matVType__3_3}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/package.scala 80:41]
  wire [127:0] ot1_tg4_matrix_b_mat_data_hi = {ot1_tg4_matrix_b_matVType__0_0,ot1_tg4_matrix_b_matVType__1_0,
    ot1_tg4_matrix_b_matVType__2_0,ot1_tg4_matrix_b_matVType__3_0,ot1_tg4_matrix_b_matVType__0_1,
    ot1_tg4_matrix_b_matVType__1_1,ot1_tg4_matrix_b_matVType__2_1,ot1_tg4_matrix_b_matVType__3_1}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/package.scala 80:41]
  wire [15:0] ot0_tg0_matrix_b_matVType_1_0_0 = io_in_bits_tc1_ot0_tg0_matrix_b[255:240]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/package.scala 77:32]
  wire [15:0] ot0_tg0_matrix_b_matVType_1_0_1 = io_in_bits_tc1_ot0_tg0_matrix_b[239:224]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/package.scala 77:32]
  wire [15:0] ot0_tg0_matrix_b_matVType_1_0_2 = io_in_bits_tc1_ot0_tg0_matrix_b[223:208]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/package.scala 77:32]
  wire [15:0] ot0_tg0_matrix_b_matVType_1_0_3 = io_in_bits_tc1_ot0_tg0_matrix_b[207:192]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/package.scala 77:32]
  wire [15:0] ot0_tg0_matrix_b_matVType_1_1_0 = io_in_bits_tc1_ot0_tg0_matrix_b[191:176]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/package.scala 77:32]
  wire [15:0] ot0_tg0_matrix_b_matVType_1_1_1 = io_in_bits_tc1_ot0_tg0_matrix_b[175:160]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/package.scala 77:32]
  wire [15:0] ot0_tg0_matrix_b_matVType_1_1_2 = io_in_bits_tc1_ot0_tg0_matrix_b[159:144]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/package.scala 77:32]
  wire [15:0] ot0_tg0_matrix_b_matVType_1_1_3 = io_in_bits_tc1_ot0_tg0_matrix_b[143:128]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/package.scala 77:32]
  wire [15:0] ot0_tg0_matrix_b_matVType_1_2_0 = io_in_bits_tc1_ot0_tg0_matrix_b[127:112]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/package.scala 77:32]
  wire [15:0] ot0_tg0_matrix_b_matVType_1_2_1 = io_in_bits_tc1_ot0_tg0_matrix_b[111:96]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/package.scala 77:32]
  wire [15:0] ot0_tg0_matrix_b_matVType_1_2_2 = io_in_bits_tc1_ot0_tg0_matrix_b[95:80]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/package.scala 77:32]
  wire [15:0] ot0_tg0_matrix_b_matVType_1_2_3 = io_in_bits_tc1_ot0_tg0_matrix_b[79:64]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/package.scala 77:32]
  wire [15:0] ot0_tg0_matrix_b_matVType_1_3_0 = io_in_bits_tc1_ot0_tg0_matrix_b[63:48]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/package.scala 77:32]
  wire [15:0] ot0_tg0_matrix_b_matVType_1_3_1 = io_in_bits_tc1_ot0_tg0_matrix_b[47:32]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/package.scala 77:32]
  wire [15:0] ot0_tg0_matrix_b_matVType_1_3_2 = io_in_bits_tc1_ot0_tg0_matrix_b[31:16]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/package.scala 77:32]
  wire [15:0] ot0_tg0_matrix_b_matVType_1_3_3 = io_in_bits_tc1_ot0_tg0_matrix_b[15:0]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/package.scala 77:32]
  wire [127:0] ot0_tg0_matrix_b_mat_data_lo_1 = {ot0_tg0_matrix_b_matVType_1_0_2,ot0_tg0_matrix_b_matVType_1_1_2,
    ot0_tg0_matrix_b_matVType_1_2_2,ot0_tg0_matrix_b_matVType_1_3_2,ot0_tg0_matrix_b_matVType_1_0_3,
    ot0_tg0_matrix_b_matVType_1_1_3,ot0_tg0_matrix_b_matVType_1_2_3,ot0_tg0_matrix_b_matVType_1_3_3}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/package.scala 80:41]
  wire [127:0] ot0_tg0_matrix_b_mat_data_hi_1 = {ot0_tg0_matrix_b_matVType_1_0_0,ot0_tg0_matrix_b_matVType_1_1_0,
    ot0_tg0_matrix_b_matVType_1_2_0,ot0_tg0_matrix_b_matVType_1_3_0,ot0_tg0_matrix_b_matVType_1_0_1,
    ot0_tg0_matrix_b_matVType_1_1_1,ot0_tg0_matrix_b_matVType_1_2_1,ot0_tg0_matrix_b_matVType_1_3_1}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/package.scala 80:41]
  wire [15:0] ot0_tg4_matrix_b_matVType_1_0_0 = io_in_bits_tc1_ot0_tg4_matrix_b[255:240]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/package.scala 77:32]
  wire [15:0] ot0_tg4_matrix_b_matVType_1_0_1 = io_in_bits_tc1_ot0_tg4_matrix_b[239:224]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/package.scala 77:32]
  wire [15:0] ot0_tg4_matrix_b_matVType_1_0_2 = io_in_bits_tc1_ot0_tg4_matrix_b[223:208]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/package.scala 77:32]
  wire [15:0] ot0_tg4_matrix_b_matVType_1_0_3 = io_in_bits_tc1_ot0_tg4_matrix_b[207:192]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/package.scala 77:32]
  wire [15:0] ot0_tg4_matrix_b_matVType_1_1_0 = io_in_bits_tc1_ot0_tg4_matrix_b[191:176]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/package.scala 77:32]
  wire [15:0] ot0_tg4_matrix_b_matVType_1_1_1 = io_in_bits_tc1_ot0_tg4_matrix_b[175:160]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/package.scala 77:32]
  wire [15:0] ot0_tg4_matrix_b_matVType_1_1_2 = io_in_bits_tc1_ot0_tg4_matrix_b[159:144]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/package.scala 77:32]
  wire [15:0] ot0_tg4_matrix_b_matVType_1_1_3 = io_in_bits_tc1_ot0_tg4_matrix_b[143:128]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/package.scala 77:32]
  wire [15:0] ot0_tg4_matrix_b_matVType_1_2_0 = io_in_bits_tc1_ot0_tg4_matrix_b[127:112]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/package.scala 77:32]
  wire [15:0] ot0_tg4_matrix_b_matVType_1_2_1 = io_in_bits_tc1_ot0_tg4_matrix_b[111:96]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/package.scala 77:32]
  wire [15:0] ot0_tg4_matrix_b_matVType_1_2_2 = io_in_bits_tc1_ot0_tg4_matrix_b[95:80]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/package.scala 77:32]
  wire [15:0] ot0_tg4_matrix_b_matVType_1_2_3 = io_in_bits_tc1_ot0_tg4_matrix_b[79:64]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/package.scala 77:32]
  wire [15:0] ot0_tg4_matrix_b_matVType_1_3_0 = io_in_bits_tc1_ot0_tg4_matrix_b[63:48]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/package.scala 77:32]
  wire [15:0] ot0_tg4_matrix_b_matVType_1_3_1 = io_in_bits_tc1_ot0_tg4_matrix_b[47:32]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/package.scala 77:32]
  wire [15:0] ot0_tg4_matrix_b_matVType_1_3_2 = io_in_bits_tc1_ot0_tg4_matrix_b[31:16]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/package.scala 77:32]
  wire [15:0] ot0_tg4_matrix_b_matVType_1_3_3 = io_in_bits_tc1_ot0_tg4_matrix_b[15:0]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/package.scala 77:32]
  wire [127:0] ot0_tg4_matrix_b_mat_data_lo_1 = {ot0_tg4_matrix_b_matVType_1_0_2,ot0_tg4_matrix_b_matVType_1_1_2,
    ot0_tg4_matrix_b_matVType_1_2_2,ot0_tg4_matrix_b_matVType_1_3_2,ot0_tg4_matrix_b_matVType_1_0_3,
    ot0_tg4_matrix_b_matVType_1_1_3,ot0_tg4_matrix_b_matVType_1_2_3,ot0_tg4_matrix_b_matVType_1_3_3}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/package.scala 80:41]
  wire [127:0] ot0_tg4_matrix_b_mat_data_hi_1 = {ot0_tg4_matrix_b_matVType_1_0_0,ot0_tg4_matrix_b_matVType_1_1_0,
    ot0_tg4_matrix_b_matVType_1_2_0,ot0_tg4_matrix_b_matVType_1_3_0,ot0_tg4_matrix_b_matVType_1_0_1,
    ot0_tg4_matrix_b_matVType_1_1_1,ot0_tg4_matrix_b_matVType_1_2_1,ot0_tg4_matrix_b_matVType_1_3_1}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/package.scala 80:41]
  wire [15:0] ot1_tg0_matrix_b_matVType_1_0_0 = io_in_bits_tc1_ot1_tg0_matrix_b[255:240]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/package.scala 77:32]
  wire [15:0] ot1_tg0_matrix_b_matVType_1_0_1 = io_in_bits_tc1_ot1_tg0_matrix_b[239:224]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/package.scala 77:32]
  wire [15:0] ot1_tg0_matrix_b_matVType_1_0_2 = io_in_bits_tc1_ot1_tg0_matrix_b[223:208]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/package.scala 77:32]
  wire [15:0] ot1_tg0_matrix_b_matVType_1_0_3 = io_in_bits_tc1_ot1_tg0_matrix_b[207:192]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/package.scala 77:32]
  wire [15:0] ot1_tg0_matrix_b_matVType_1_1_0 = io_in_bits_tc1_ot1_tg0_matrix_b[191:176]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/package.scala 77:32]
  wire [15:0] ot1_tg0_matrix_b_matVType_1_1_1 = io_in_bits_tc1_ot1_tg0_matrix_b[175:160]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/package.scala 77:32]
  wire [15:0] ot1_tg0_matrix_b_matVType_1_1_2 = io_in_bits_tc1_ot1_tg0_matrix_b[159:144]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/package.scala 77:32]
  wire [15:0] ot1_tg0_matrix_b_matVType_1_1_3 = io_in_bits_tc1_ot1_tg0_matrix_b[143:128]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/package.scala 77:32]
  wire [15:0] ot1_tg0_matrix_b_matVType_1_2_0 = io_in_bits_tc1_ot1_tg0_matrix_b[127:112]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/package.scala 77:32]
  wire [15:0] ot1_tg0_matrix_b_matVType_1_2_1 = io_in_bits_tc1_ot1_tg0_matrix_b[111:96]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/package.scala 77:32]
  wire [15:0] ot1_tg0_matrix_b_matVType_1_2_2 = io_in_bits_tc1_ot1_tg0_matrix_b[95:80]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/package.scala 77:32]
  wire [15:0] ot1_tg0_matrix_b_matVType_1_2_3 = io_in_bits_tc1_ot1_tg0_matrix_b[79:64]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/package.scala 77:32]
  wire [15:0] ot1_tg0_matrix_b_matVType_1_3_0 = io_in_bits_tc1_ot1_tg0_matrix_b[63:48]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/package.scala 77:32]
  wire [15:0] ot1_tg0_matrix_b_matVType_1_3_1 = io_in_bits_tc1_ot1_tg0_matrix_b[47:32]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/package.scala 77:32]
  wire [15:0] ot1_tg0_matrix_b_matVType_1_3_2 = io_in_bits_tc1_ot1_tg0_matrix_b[31:16]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/package.scala 77:32]
  wire [15:0] ot1_tg0_matrix_b_matVType_1_3_3 = io_in_bits_tc1_ot1_tg0_matrix_b[15:0]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/package.scala 77:32]
  wire [127:0] ot1_tg0_matrix_b_mat_data_lo_1 = {ot1_tg0_matrix_b_matVType_1_0_2,ot1_tg0_matrix_b_matVType_1_1_2,
    ot1_tg0_matrix_b_matVType_1_2_2,ot1_tg0_matrix_b_matVType_1_3_2,ot1_tg0_matrix_b_matVType_1_0_3,
    ot1_tg0_matrix_b_matVType_1_1_3,ot1_tg0_matrix_b_matVType_1_2_3,ot1_tg0_matrix_b_matVType_1_3_3}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/package.scala 80:41]
  wire [127:0] ot1_tg0_matrix_b_mat_data_hi_1 = {ot1_tg0_matrix_b_matVType_1_0_0,ot1_tg0_matrix_b_matVType_1_1_0,
    ot1_tg0_matrix_b_matVType_1_2_0,ot1_tg0_matrix_b_matVType_1_3_0,ot1_tg0_matrix_b_matVType_1_0_1,
    ot1_tg0_matrix_b_matVType_1_1_1,ot1_tg0_matrix_b_matVType_1_2_1,ot1_tg0_matrix_b_matVType_1_3_1}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/package.scala 80:41]
  wire [15:0] ot1_tg4_matrix_b_matVType_1_0_0 = io_in_bits_tc1_ot1_tg4_matrix_b[255:240]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/package.scala 77:32]
  wire [15:0] ot1_tg4_matrix_b_matVType_1_0_1 = io_in_bits_tc1_ot1_tg4_matrix_b[239:224]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/package.scala 77:32]
  wire [15:0] ot1_tg4_matrix_b_matVType_1_0_2 = io_in_bits_tc1_ot1_tg4_matrix_b[223:208]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/package.scala 77:32]
  wire [15:0] ot1_tg4_matrix_b_matVType_1_0_3 = io_in_bits_tc1_ot1_tg4_matrix_b[207:192]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/package.scala 77:32]
  wire [15:0] ot1_tg4_matrix_b_matVType_1_1_0 = io_in_bits_tc1_ot1_tg4_matrix_b[191:176]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/package.scala 77:32]
  wire [15:0] ot1_tg4_matrix_b_matVType_1_1_1 = io_in_bits_tc1_ot1_tg4_matrix_b[175:160]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/package.scala 77:32]
  wire [15:0] ot1_tg4_matrix_b_matVType_1_1_2 = io_in_bits_tc1_ot1_tg4_matrix_b[159:144]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/package.scala 77:32]
  wire [15:0] ot1_tg4_matrix_b_matVType_1_1_3 = io_in_bits_tc1_ot1_tg4_matrix_b[143:128]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/package.scala 77:32]
  wire [15:0] ot1_tg4_matrix_b_matVType_1_2_0 = io_in_bits_tc1_ot1_tg4_matrix_b[127:112]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/package.scala 77:32]
  wire [15:0] ot1_tg4_matrix_b_matVType_1_2_1 = io_in_bits_tc1_ot1_tg4_matrix_b[111:96]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/package.scala 77:32]
  wire [15:0] ot1_tg4_matrix_b_matVType_1_2_2 = io_in_bits_tc1_ot1_tg4_matrix_b[95:80]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/package.scala 77:32]
  wire [15:0] ot1_tg4_matrix_b_matVType_1_2_3 = io_in_bits_tc1_ot1_tg4_matrix_b[79:64]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/package.scala 77:32]
  wire [15:0] ot1_tg4_matrix_b_matVType_1_3_0 = io_in_bits_tc1_ot1_tg4_matrix_b[63:48]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/package.scala 77:32]
  wire [15:0] ot1_tg4_matrix_b_matVType_1_3_1 = io_in_bits_tc1_ot1_tg4_matrix_b[47:32]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/package.scala 77:32]
  wire [15:0] ot1_tg4_matrix_b_matVType_1_3_2 = io_in_bits_tc1_ot1_tg4_matrix_b[31:16]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/package.scala 77:32]
  wire [15:0] ot1_tg4_matrix_b_matVType_1_3_3 = io_in_bits_tc1_ot1_tg4_matrix_b[15:0]; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/package.scala 77:32]
  wire [127:0] ot1_tg4_matrix_b_mat_data_lo_1 = {ot1_tg4_matrix_b_matVType_1_0_2,ot1_tg4_matrix_b_matVType_1_1_2,
    ot1_tg4_matrix_b_matVType_1_2_2,ot1_tg4_matrix_b_matVType_1_3_2,ot1_tg4_matrix_b_matVType_1_0_3,
    ot1_tg4_matrix_b_matVType_1_1_3,ot1_tg4_matrix_b_matVType_1_2_3,ot1_tg4_matrix_b_matVType_1_3_3}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/package.scala 80:41]
  wire [127:0] ot1_tg4_matrix_b_mat_data_hi_1 = {ot1_tg4_matrix_b_matVType_1_0_0,ot1_tg4_matrix_b_matVType_1_1_0,
    ot1_tg4_matrix_b_matVType_1_2_0,ot1_tg4_matrix_b_matVType_1_3_0,ot1_tg4_matrix_b_matVType_1_0_1,
    ot1_tg4_matrix_b_matVType_1_1_1,ot1_tg4_matrix_b_matVType_1_2_1,ot1_tg4_matrix_b_matVType_1_3_1}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/package.scala 80:41]
  wire  tc_ready_0 = tc_io_in_ready; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/Top.scala 59:22 86:17]
  wire  tc_ready_1 = tc_1_io_in_ready; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/Top.scala 59:22 86:17]
  wire  tc_valid_0 = tc_io_out_valid; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/Top.scala 58:22 85:17]
  wire  tc_valid_1 = tc_1_io_out_valid; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/Top.scala 58:22 85:17]
  TensorCore tc ( // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/TensorCore.scala 67:20]
    .clock(tc_clock),
    .reset(tc_reset),
    .io_in_ready(tc_io_in_ready),
    .io_in_valid(tc_io_in_valid),
    .io_in_bits_octet0_threadgroup0_matrix_a_data(tc_io_in_bits_octet0_threadgroup0_matrix_a_data),
    .io_in_bits_octet0_threadgroup0_matrix_b_data(tc_io_in_bits_octet0_threadgroup0_matrix_b_data),
    .io_in_bits_octet0_threadgroup0_matrix_c_data(tc_io_in_bits_octet0_threadgroup0_matrix_c_data),
    .io_in_bits_octet0_threadgroup4_matrix_a_data(tc_io_in_bits_octet0_threadgroup4_matrix_a_data),
    .io_in_bits_octet0_threadgroup4_matrix_b_data(tc_io_in_bits_octet0_threadgroup4_matrix_b_data),
    .io_in_bits_octet0_threadgroup4_matrix_c_data(tc_io_in_bits_octet0_threadgroup4_matrix_c_data),
    .io_in_bits_octet1_threadgroup0_matrix_a_data(tc_io_in_bits_octet1_threadgroup0_matrix_a_data),
    .io_in_bits_octet1_threadgroup0_matrix_b_data(tc_io_in_bits_octet1_threadgroup0_matrix_b_data),
    .io_in_bits_octet1_threadgroup0_matrix_c_data(tc_io_in_bits_octet1_threadgroup0_matrix_c_data),
    .io_in_bits_octet1_threadgroup4_matrix_a_data(tc_io_in_bits_octet1_threadgroup4_matrix_a_data),
    .io_in_bits_octet1_threadgroup4_matrix_b_data(tc_io_in_bits_octet1_threadgroup4_matrix_b_data),
    .io_in_bits_octet1_threadgroup4_matrix_c_data(tc_io_in_bits_octet1_threadgroup4_matrix_c_data),
    .io_in_bits_ctrl_matBSel(tc_io_in_bits_ctrl_matBSel),
    .io_in_bits_ctrl_mixPcMode(tc_io_in_bits_ctrl_mixPcMode),
    .io_out_valid(tc_io_out_valid),
    .io_out_bits_octet0_threadgroup0_matrix_d_data(tc_io_out_bits_octet0_threadgroup0_matrix_d_data),
    .io_out_bits_octet0_threadgroup4_matrix_d_data(tc_io_out_bits_octet0_threadgroup4_matrix_d_data),
    .io_out_bits_octet1_threadgroup0_matrix_d_data(tc_io_out_bits_octet1_threadgroup0_matrix_d_data),
    .io_out_bits_octet1_threadgroup4_matrix_d_data(tc_io_out_bits_octet1_threadgroup4_matrix_d_data)
  );
  TensorCore tc_1 ( // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/TensorCore.scala 67:20]
    .clock(tc_1_clock),
    .reset(tc_1_reset),
    .io_in_ready(tc_1_io_in_ready),
    .io_in_valid(tc_1_io_in_valid),
    .io_in_bits_octet0_threadgroup0_matrix_a_data(tc_1_io_in_bits_octet0_threadgroup0_matrix_a_data),
    .io_in_bits_octet0_threadgroup0_matrix_b_data(tc_1_io_in_bits_octet0_threadgroup0_matrix_b_data),
    .io_in_bits_octet0_threadgroup0_matrix_c_data(tc_1_io_in_bits_octet0_threadgroup0_matrix_c_data),
    .io_in_bits_octet0_threadgroup4_matrix_a_data(tc_1_io_in_bits_octet0_threadgroup4_matrix_a_data),
    .io_in_bits_octet0_threadgroup4_matrix_b_data(tc_1_io_in_bits_octet0_threadgroup4_matrix_b_data),
    .io_in_bits_octet0_threadgroup4_matrix_c_data(tc_1_io_in_bits_octet0_threadgroup4_matrix_c_data),
    .io_in_bits_octet1_threadgroup0_matrix_a_data(tc_1_io_in_bits_octet1_threadgroup0_matrix_a_data),
    .io_in_bits_octet1_threadgroup0_matrix_b_data(tc_1_io_in_bits_octet1_threadgroup0_matrix_b_data),
    .io_in_bits_octet1_threadgroup0_matrix_c_data(tc_1_io_in_bits_octet1_threadgroup0_matrix_c_data),
    .io_in_bits_octet1_threadgroup4_matrix_a_data(tc_1_io_in_bits_octet1_threadgroup4_matrix_a_data),
    .io_in_bits_octet1_threadgroup4_matrix_b_data(tc_1_io_in_bits_octet1_threadgroup4_matrix_b_data),
    .io_in_bits_octet1_threadgroup4_matrix_c_data(tc_1_io_in_bits_octet1_threadgroup4_matrix_c_data),
    .io_in_bits_ctrl_matBSel(tc_1_io_in_bits_ctrl_matBSel),
    .io_in_bits_ctrl_mixPcMode(tc_1_io_in_bits_ctrl_mixPcMode),
    .io_out_valid(tc_1_io_out_valid),
    .io_out_bits_octet0_threadgroup0_matrix_d_data(tc_1_io_out_bits_octet0_threadgroup0_matrix_d_data),
    .io_out_bits_octet0_threadgroup4_matrix_d_data(tc_1_io_out_bits_octet0_threadgroup4_matrix_d_data),
    .io_out_bits_octet1_threadgroup0_matrix_d_data(tc_1_io_out_bits_octet1_threadgroup0_matrix_d_data),
    .io_out_bits_octet1_threadgroup4_matrix_d_data(tc_1_io_out_bits_octet1_threadgroup4_matrix_d_data)
  );
  assign io_in_ready = tc_ready_0 & tc_ready_1; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/Top.scala 89:36]
  assign io_out_valid = tc_valid_0 & tc_valid_1; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/Top.scala 90:36]
  assign io_out_bits_tc0_octet0_threadgroup0_matrix_d_data = tc_io_out_bits_octet0_threadgroup0_matrix_d_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/Top.scala 83:{31,31}]
  assign io_out_bits_tc0_octet0_threadgroup4_matrix_d_data = tc_io_out_bits_octet0_threadgroup4_matrix_d_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/Top.scala 83:{31,31}]
  assign io_out_bits_tc0_octet1_threadgroup0_matrix_d_data = tc_io_out_bits_octet1_threadgroup0_matrix_d_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/Top.scala 84:{31,31}]
  assign io_out_bits_tc0_octet1_threadgroup4_matrix_d_data = tc_io_out_bits_octet1_threadgroup4_matrix_d_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/Top.scala 84:{31,31}]
  assign io_out_bits_tc1_octet0_threadgroup0_matrix_d_data = tc_1_io_out_bits_octet0_threadgroup0_matrix_d_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/Top.scala 83:{31,31}]
  assign io_out_bits_tc1_octet0_threadgroup4_matrix_d_data = tc_1_io_out_bits_octet0_threadgroup4_matrix_d_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/Top.scala 83:{31,31}]
  assign io_out_bits_tc1_octet1_threadgroup0_matrix_d_data = tc_1_io_out_bits_octet1_threadgroup0_matrix_d_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/Top.scala 84:{31,31}]
  assign io_out_bits_tc1_octet1_threadgroup4_matrix_d_data = tc_1_io_out_bits_octet1_threadgroup4_matrix_d_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/Top.scala 84:{31,31}]
  assign tc_clock = clock;
  assign tc_reset = reset;
  assign tc_io_in_valid = io_in_valid; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/TensorCore.scala 78:20]
  assign tc_io_in_bits_octet0_threadgroup0_matrix_a_data = io_in_bits_tc0_ot0_tg0_matrix_a; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/Top.scala 54:{27,27}]
  assign tc_io_in_bits_octet0_threadgroup0_matrix_b_data = {ot0_tg0_matrix_b_mat_data_hi,ot0_tg0_matrix_b_mat_data_lo}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/package.scala 80:41]
  assign tc_io_in_bits_octet0_threadgroup0_matrix_c_data = io_in_bits_tc0_ot0_tg0_matrix_c; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/Top.scala 54:{27,27}]
  assign tc_io_in_bits_octet0_threadgroup4_matrix_a_data = io_in_bits_tc0_ot0_tg4_matrix_a; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/Top.scala 54:{27,27}]
  assign tc_io_in_bits_octet0_threadgroup4_matrix_b_data = {ot0_tg4_matrix_b_mat_data_hi,ot0_tg4_matrix_b_mat_data_lo}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/package.scala 80:41]
  assign tc_io_in_bits_octet0_threadgroup4_matrix_c_data = io_in_bits_tc0_ot0_tg4_matrix_c; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/Top.scala 54:{27,27}]
  assign tc_io_in_bits_octet1_threadgroup0_matrix_a_data = io_in_bits_tc0_ot1_tg0_matrix_a; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/Top.scala 54:{27,27}]
  assign tc_io_in_bits_octet1_threadgroup0_matrix_b_data = {ot1_tg0_matrix_b_mat_data_hi,ot1_tg0_matrix_b_mat_data_lo}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/package.scala 80:41]
  assign tc_io_in_bits_octet1_threadgroup0_matrix_c_data = io_in_bits_tc0_ot1_tg0_matrix_c; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/Top.scala 54:{27,27}]
  assign tc_io_in_bits_octet1_threadgroup4_matrix_a_data = io_in_bits_tc0_ot1_tg4_matrix_a; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/Top.scala 54:{27,27}]
  assign tc_io_in_bits_octet1_threadgroup4_matrix_b_data = {ot1_tg4_matrix_b_mat_data_hi,ot1_tg4_matrix_b_mat_data_lo}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/package.scala 80:41]
  assign tc_io_in_bits_octet1_threadgroup4_matrix_c_data = io_in_bits_tc0_ot1_tg4_matrix_c; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/Top.scala 54:{27,27}]
  assign tc_io_in_bits_ctrl_matBSel = io_in_bits_ctrl_matBSel; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/TensorCore.scala 94:32]
  assign tc_io_in_bits_ctrl_mixPcMode = io_in_bits_ctrl_mixPcMode; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/TensorCore.scala 95:34]
  assign tc_1_clock = clock;
  assign tc_1_reset = reset;
  assign tc_1_io_in_valid = io_in_valid; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/TensorCore.scala 78:20]
  assign tc_1_io_in_bits_octet0_threadgroup0_matrix_a_data = io_in_bits_tc1_ot0_tg0_matrix_a; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/Top.scala 54:{27,27}]
  assign tc_1_io_in_bits_octet0_threadgroup0_matrix_b_data = {ot0_tg0_matrix_b_mat_data_hi_1,
    ot0_tg0_matrix_b_mat_data_lo_1}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/package.scala 80:41]
  assign tc_1_io_in_bits_octet0_threadgroup0_matrix_c_data = io_in_bits_tc1_ot0_tg0_matrix_c; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/Top.scala 54:{27,27}]
  assign tc_1_io_in_bits_octet0_threadgroup4_matrix_a_data = io_in_bits_tc1_ot0_tg4_matrix_a; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/Top.scala 54:{27,27}]
  assign tc_1_io_in_bits_octet0_threadgroup4_matrix_b_data = {ot0_tg4_matrix_b_mat_data_hi_1,
    ot0_tg4_matrix_b_mat_data_lo_1}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/package.scala 80:41]
  assign tc_1_io_in_bits_octet0_threadgroup4_matrix_c_data = io_in_bits_tc1_ot0_tg4_matrix_c; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/Top.scala 54:{27,27}]
  assign tc_1_io_in_bits_octet1_threadgroup0_matrix_a_data = io_in_bits_tc1_ot1_tg0_matrix_a; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/Top.scala 54:{27,27}]
  assign tc_1_io_in_bits_octet1_threadgroup0_matrix_b_data = {ot1_tg0_matrix_b_mat_data_hi_1,
    ot1_tg0_matrix_b_mat_data_lo_1}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/package.scala 80:41]
  assign tc_1_io_in_bits_octet1_threadgroup0_matrix_c_data = io_in_bits_tc1_ot1_tg0_matrix_c; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/Top.scala 54:{27,27}]
  assign tc_1_io_in_bits_octet1_threadgroup4_matrix_a_data = io_in_bits_tc1_ot1_tg4_matrix_a; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/Top.scala 54:{27,27}]
  assign tc_1_io_in_bits_octet1_threadgroup4_matrix_b_data = {ot1_tg4_matrix_b_mat_data_hi_1,
    ot1_tg4_matrix_b_mat_data_lo_1}; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/package.scala 80:41]
  assign tc_1_io_in_bits_octet1_threadgroup4_matrix_c_data = io_in_bits_tc1_ot1_tg4_matrix_c; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/Top.scala 54:{27,27}]
  assign tc_1_io_in_bits_ctrl_matBSel = io_in_bits_ctrl_matBSel; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/TensorCore.scala 94:32]
  assign tc_1_io_in_bits_ctrl_mixPcMode = io_in_bits_ctrl_mixPcMode; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/TensorCore/TensorCore.scala 95:34]
endmodule
module Adagio(
  input         clock,
  input         reset,
  input         io_mixPc, // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Adagio.scala 11:14]
  input         io_uart_ctrl_tx_done, // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Adagio.scala 11:14]
  input         io_uart_ctrl_rx_valid, // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Adagio.scala 11:14]
  output        io_uart_ctrl_tx_en, // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Adagio.scala 11:14]
  input         io_rf_w_en, // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Adagio.scala 11:14]
  input  [7:0]  io_rf_r_addr, // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Adagio.scala 11:14]
  input  [7:0]  io_rf_w_addr, // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Adagio.scala 11:14]
  output [63:0] io_rf_r_data, // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Adagio.scala 11:14]
  input  [63:0] io_rf_w_data // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Adagio.scala 11:14]
);
  wire  manager_clock; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Adagio.scala 16:23]
  wire  manager_reset; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Adagio.scala 16:23]
  wire  manager_io_mixPc; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Adagio.scala 16:23]
  wire  manager_io_uart_ctrl_tx_done; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Adagio.scala 16:23]
  wire  manager_io_uart_ctrl_rx_valid; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Adagio.scala 16:23]
  wire  manager_io_uart_ctrl_tx_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Adagio.scala 16:23]
  wire  manager_io_uart_rf_w_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Adagio.scala 16:23]
  wire [7:0] manager_io_uart_rf_r_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Adagio.scala 16:23]
  wire [7:0] manager_io_uart_rf_w_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Adagio.scala 16:23]
  wire [63:0] manager_io_uart_rf_r_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Adagio.scala 16:23]
  wire [63:0] manager_io_uart_rf_w_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Adagio.scala 16:23]
  wire  manager_io_top_src_ready; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Adagio.scala 16:23]
  wire  manager_io_top_src_valid; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Adagio.scala 16:23]
  wire [255:0] manager_io_top_src_bits_tc0_ot0_tg0_matrix_a; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Adagio.scala 16:23]
  wire [255:0] manager_io_top_src_bits_tc0_ot0_tg0_matrix_b; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Adagio.scala 16:23]
  wire [255:0] manager_io_top_src_bits_tc0_ot0_tg0_matrix_c; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Adagio.scala 16:23]
  wire [255:0] manager_io_top_src_bits_tc0_ot0_tg4_matrix_a; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Adagio.scala 16:23]
  wire [255:0] manager_io_top_src_bits_tc0_ot0_tg4_matrix_b; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Adagio.scala 16:23]
  wire [255:0] manager_io_top_src_bits_tc0_ot0_tg4_matrix_c; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Adagio.scala 16:23]
  wire [255:0] manager_io_top_src_bits_tc0_ot1_tg0_matrix_a; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Adagio.scala 16:23]
  wire [255:0] manager_io_top_src_bits_tc0_ot1_tg0_matrix_b; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Adagio.scala 16:23]
  wire [255:0] manager_io_top_src_bits_tc0_ot1_tg0_matrix_c; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Adagio.scala 16:23]
  wire [255:0] manager_io_top_src_bits_tc0_ot1_tg4_matrix_a; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Adagio.scala 16:23]
  wire [255:0] manager_io_top_src_bits_tc0_ot1_tg4_matrix_b; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Adagio.scala 16:23]
  wire [255:0] manager_io_top_src_bits_tc0_ot1_tg4_matrix_c; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Adagio.scala 16:23]
  wire [255:0] manager_io_top_src_bits_tc1_ot0_tg0_matrix_a; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Adagio.scala 16:23]
  wire [255:0] manager_io_top_src_bits_tc1_ot0_tg0_matrix_b; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Adagio.scala 16:23]
  wire [255:0] manager_io_top_src_bits_tc1_ot0_tg0_matrix_c; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Adagio.scala 16:23]
  wire [255:0] manager_io_top_src_bits_tc1_ot0_tg4_matrix_a; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Adagio.scala 16:23]
  wire [255:0] manager_io_top_src_bits_tc1_ot0_tg4_matrix_b; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Adagio.scala 16:23]
  wire [255:0] manager_io_top_src_bits_tc1_ot0_tg4_matrix_c; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Adagio.scala 16:23]
  wire [255:0] manager_io_top_src_bits_tc1_ot1_tg0_matrix_a; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Adagio.scala 16:23]
  wire [255:0] manager_io_top_src_bits_tc1_ot1_tg0_matrix_b; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Adagio.scala 16:23]
  wire [255:0] manager_io_top_src_bits_tc1_ot1_tg0_matrix_c; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Adagio.scala 16:23]
  wire [255:0] manager_io_top_src_bits_tc1_ot1_tg4_matrix_a; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Adagio.scala 16:23]
  wire [255:0] manager_io_top_src_bits_tc1_ot1_tg4_matrix_b; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Adagio.scala 16:23]
  wire [255:0] manager_io_top_src_bits_tc1_ot1_tg4_matrix_c; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Adagio.scala 16:23]
  wire  manager_io_top_src_bits_ctrl_matBSel; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Adagio.scala 16:23]
  wire  manager_io_top_src_bits_ctrl_mixPcMode; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Adagio.scala 16:23]
  wire  manager_io_top_wb_ready; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Adagio.scala 16:23]
  wire  manager_io_top_wb_valid; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Adagio.scala 16:23]
  wire [255:0] manager_io_top_wb_bits_tc0_octet0_threadgroup0_matrix_d_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Adagio.scala 16:23]
  wire [255:0] manager_io_top_wb_bits_tc0_octet0_threadgroup4_matrix_d_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Adagio.scala 16:23]
  wire [255:0] manager_io_top_wb_bits_tc0_octet1_threadgroup0_matrix_d_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Adagio.scala 16:23]
  wire [255:0] manager_io_top_wb_bits_tc0_octet1_threadgroup4_matrix_d_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Adagio.scala 16:23]
  wire [255:0] manager_io_top_wb_bits_tc1_octet0_threadgroup0_matrix_d_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Adagio.scala 16:23]
  wire [255:0] manager_io_top_wb_bits_tc1_octet0_threadgroup4_matrix_d_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Adagio.scala 16:23]
  wire [255:0] manager_io_top_wb_bits_tc1_octet1_threadgroup0_matrix_d_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Adagio.scala 16:23]
  wire [255:0] manager_io_top_wb_bits_tc1_octet1_threadgroup4_matrix_d_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Adagio.scala 16:23]
  wire  top_clock; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Adagio.scala 17:19]
  wire  top_reset; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Adagio.scala 17:19]
  wire  top_io_in_ready; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Adagio.scala 17:19]
  wire  top_io_in_valid; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Adagio.scala 17:19]
  wire [255:0] top_io_in_bits_tc0_ot0_tg0_matrix_a; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Adagio.scala 17:19]
  wire [255:0] top_io_in_bits_tc0_ot0_tg0_matrix_b; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Adagio.scala 17:19]
  wire [255:0] top_io_in_bits_tc0_ot0_tg0_matrix_c; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Adagio.scala 17:19]
  wire [255:0] top_io_in_bits_tc0_ot0_tg4_matrix_a; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Adagio.scala 17:19]
  wire [255:0] top_io_in_bits_tc0_ot0_tg4_matrix_b; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Adagio.scala 17:19]
  wire [255:0] top_io_in_bits_tc0_ot0_tg4_matrix_c; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Adagio.scala 17:19]
  wire [255:0] top_io_in_bits_tc0_ot1_tg0_matrix_a; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Adagio.scala 17:19]
  wire [255:0] top_io_in_bits_tc0_ot1_tg0_matrix_b; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Adagio.scala 17:19]
  wire [255:0] top_io_in_bits_tc0_ot1_tg0_matrix_c; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Adagio.scala 17:19]
  wire [255:0] top_io_in_bits_tc0_ot1_tg4_matrix_a; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Adagio.scala 17:19]
  wire [255:0] top_io_in_bits_tc0_ot1_tg4_matrix_b; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Adagio.scala 17:19]
  wire [255:0] top_io_in_bits_tc0_ot1_tg4_matrix_c; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Adagio.scala 17:19]
  wire [255:0] top_io_in_bits_tc1_ot0_tg0_matrix_a; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Adagio.scala 17:19]
  wire [255:0] top_io_in_bits_tc1_ot0_tg0_matrix_b; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Adagio.scala 17:19]
  wire [255:0] top_io_in_bits_tc1_ot0_tg0_matrix_c; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Adagio.scala 17:19]
  wire [255:0] top_io_in_bits_tc1_ot0_tg4_matrix_a; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Adagio.scala 17:19]
  wire [255:0] top_io_in_bits_tc1_ot0_tg4_matrix_b; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Adagio.scala 17:19]
  wire [255:0] top_io_in_bits_tc1_ot0_tg4_matrix_c; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Adagio.scala 17:19]
  wire [255:0] top_io_in_bits_tc1_ot1_tg0_matrix_a; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Adagio.scala 17:19]
  wire [255:0] top_io_in_bits_tc1_ot1_tg0_matrix_b; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Adagio.scala 17:19]
  wire [255:0] top_io_in_bits_tc1_ot1_tg0_matrix_c; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Adagio.scala 17:19]
  wire [255:0] top_io_in_bits_tc1_ot1_tg4_matrix_a; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Adagio.scala 17:19]
  wire [255:0] top_io_in_bits_tc1_ot1_tg4_matrix_b; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Adagio.scala 17:19]
  wire [255:0] top_io_in_bits_tc1_ot1_tg4_matrix_c; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Adagio.scala 17:19]
  wire  top_io_in_bits_ctrl_matBSel; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Adagio.scala 17:19]
  wire  top_io_in_bits_ctrl_mixPcMode; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Adagio.scala 17:19]
  wire  top_io_out_valid; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Adagio.scala 17:19]
  wire [255:0] top_io_out_bits_tc0_octet0_threadgroup0_matrix_d_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Adagio.scala 17:19]
  wire [255:0] top_io_out_bits_tc0_octet0_threadgroup4_matrix_d_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Adagio.scala 17:19]
  wire [255:0] top_io_out_bits_tc0_octet1_threadgroup0_matrix_d_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Adagio.scala 17:19]
  wire [255:0] top_io_out_bits_tc0_octet1_threadgroup4_matrix_d_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Adagio.scala 17:19]
  wire [255:0] top_io_out_bits_tc1_octet0_threadgroup0_matrix_d_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Adagio.scala 17:19]
  wire [255:0] top_io_out_bits_tc1_octet0_threadgroup4_matrix_d_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Adagio.scala 17:19]
  wire [255:0] top_io_out_bits_tc1_octet1_threadgroup0_matrix_d_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Adagio.scala 17:19]
  wire [255:0] top_io_out_bits_tc1_octet1_threadgroup4_matrix_d_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Adagio.scala 17:19]
  Manager manager ( // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Adagio.scala 16:23]
    .clock(manager_clock),
    .reset(manager_reset),
    .io_mixPc(manager_io_mixPc),
    .io_uart_ctrl_tx_done(manager_io_uart_ctrl_tx_done),
    .io_uart_ctrl_rx_valid(manager_io_uart_ctrl_rx_valid),
    .io_uart_ctrl_tx_en(manager_io_uart_ctrl_tx_en),
    .io_uart_rf_w_en(manager_io_uart_rf_w_en),
    .io_uart_rf_r_addr(manager_io_uart_rf_r_addr),
    .io_uart_rf_w_addr(manager_io_uart_rf_w_addr),
    .io_uart_rf_r_data(manager_io_uart_rf_r_data),
    .io_uart_rf_w_data(manager_io_uart_rf_w_data),
    .io_top_src_ready(manager_io_top_src_ready),
    .io_top_src_valid(manager_io_top_src_valid),
    .io_top_src_bits_tc0_ot0_tg0_matrix_a(manager_io_top_src_bits_tc0_ot0_tg0_matrix_a),
    .io_top_src_bits_tc0_ot0_tg0_matrix_b(manager_io_top_src_bits_tc0_ot0_tg0_matrix_b),
    .io_top_src_bits_tc0_ot0_tg0_matrix_c(manager_io_top_src_bits_tc0_ot0_tg0_matrix_c),
    .io_top_src_bits_tc0_ot0_tg4_matrix_a(manager_io_top_src_bits_tc0_ot0_tg4_matrix_a),
    .io_top_src_bits_tc0_ot0_tg4_matrix_b(manager_io_top_src_bits_tc0_ot0_tg4_matrix_b),
    .io_top_src_bits_tc0_ot0_tg4_matrix_c(manager_io_top_src_bits_tc0_ot0_tg4_matrix_c),
    .io_top_src_bits_tc0_ot1_tg0_matrix_a(manager_io_top_src_bits_tc0_ot1_tg0_matrix_a),
    .io_top_src_bits_tc0_ot1_tg0_matrix_b(manager_io_top_src_bits_tc0_ot1_tg0_matrix_b),
    .io_top_src_bits_tc0_ot1_tg0_matrix_c(manager_io_top_src_bits_tc0_ot1_tg0_matrix_c),
    .io_top_src_bits_tc0_ot1_tg4_matrix_a(manager_io_top_src_bits_tc0_ot1_tg4_matrix_a),
    .io_top_src_bits_tc0_ot1_tg4_matrix_b(manager_io_top_src_bits_tc0_ot1_tg4_matrix_b),
    .io_top_src_bits_tc0_ot1_tg4_matrix_c(manager_io_top_src_bits_tc0_ot1_tg4_matrix_c),
    .io_top_src_bits_tc1_ot0_tg0_matrix_a(manager_io_top_src_bits_tc1_ot0_tg0_matrix_a),
    .io_top_src_bits_tc1_ot0_tg0_matrix_b(manager_io_top_src_bits_tc1_ot0_tg0_matrix_b),
    .io_top_src_bits_tc1_ot0_tg0_matrix_c(manager_io_top_src_bits_tc1_ot0_tg0_matrix_c),
    .io_top_src_bits_tc1_ot0_tg4_matrix_a(manager_io_top_src_bits_tc1_ot0_tg4_matrix_a),
    .io_top_src_bits_tc1_ot0_tg4_matrix_b(manager_io_top_src_bits_tc1_ot0_tg4_matrix_b),
    .io_top_src_bits_tc1_ot0_tg4_matrix_c(manager_io_top_src_bits_tc1_ot0_tg4_matrix_c),
    .io_top_src_bits_tc1_ot1_tg0_matrix_a(manager_io_top_src_bits_tc1_ot1_tg0_matrix_a),
    .io_top_src_bits_tc1_ot1_tg0_matrix_b(manager_io_top_src_bits_tc1_ot1_tg0_matrix_b),
    .io_top_src_bits_tc1_ot1_tg0_matrix_c(manager_io_top_src_bits_tc1_ot1_tg0_matrix_c),
    .io_top_src_bits_tc1_ot1_tg4_matrix_a(manager_io_top_src_bits_tc1_ot1_tg4_matrix_a),
    .io_top_src_bits_tc1_ot1_tg4_matrix_b(manager_io_top_src_bits_tc1_ot1_tg4_matrix_b),
    .io_top_src_bits_tc1_ot1_tg4_matrix_c(manager_io_top_src_bits_tc1_ot1_tg4_matrix_c),
    .io_top_src_bits_ctrl_matBSel(manager_io_top_src_bits_ctrl_matBSel),
    .io_top_src_bits_ctrl_mixPcMode(manager_io_top_src_bits_ctrl_mixPcMode),
    .io_top_wb_ready(manager_io_top_wb_ready),
    .io_top_wb_valid(manager_io_top_wb_valid),
    .io_top_wb_bits_tc0_octet0_threadgroup0_matrix_d_data(manager_io_top_wb_bits_tc0_octet0_threadgroup0_matrix_d_data),
    .io_top_wb_bits_tc0_octet0_threadgroup4_matrix_d_data(manager_io_top_wb_bits_tc0_octet0_threadgroup4_matrix_d_data),
    .io_top_wb_bits_tc0_octet1_threadgroup0_matrix_d_data(manager_io_top_wb_bits_tc0_octet1_threadgroup0_matrix_d_data),
    .io_top_wb_bits_tc0_octet1_threadgroup4_matrix_d_data(manager_io_top_wb_bits_tc0_octet1_threadgroup4_matrix_d_data),
    .io_top_wb_bits_tc1_octet0_threadgroup0_matrix_d_data(manager_io_top_wb_bits_tc1_octet0_threadgroup0_matrix_d_data),
    .io_top_wb_bits_tc1_octet0_threadgroup4_matrix_d_data(manager_io_top_wb_bits_tc1_octet0_threadgroup4_matrix_d_data),
    .io_top_wb_bits_tc1_octet1_threadgroup0_matrix_d_data(manager_io_top_wb_bits_tc1_octet1_threadgroup0_matrix_d_data),
    .io_top_wb_bits_tc1_octet1_threadgroup4_matrix_d_data(manager_io_top_wb_bits_tc1_octet1_threadgroup4_matrix_d_data)
  );
  Top top ( // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Adagio.scala 17:19]
    .clock(top_clock),
    .reset(top_reset),
    .io_in_ready(top_io_in_ready),
    .io_in_valid(top_io_in_valid),
    .io_in_bits_tc0_ot0_tg0_matrix_a(top_io_in_bits_tc0_ot0_tg0_matrix_a),
    .io_in_bits_tc0_ot0_tg0_matrix_b(top_io_in_bits_tc0_ot0_tg0_matrix_b),
    .io_in_bits_tc0_ot0_tg0_matrix_c(top_io_in_bits_tc0_ot0_tg0_matrix_c),
    .io_in_bits_tc0_ot0_tg4_matrix_a(top_io_in_bits_tc0_ot0_tg4_matrix_a),
    .io_in_bits_tc0_ot0_tg4_matrix_b(top_io_in_bits_tc0_ot0_tg4_matrix_b),
    .io_in_bits_tc0_ot0_tg4_matrix_c(top_io_in_bits_tc0_ot0_tg4_matrix_c),
    .io_in_bits_tc0_ot1_tg0_matrix_a(top_io_in_bits_tc0_ot1_tg0_matrix_a),
    .io_in_bits_tc0_ot1_tg0_matrix_b(top_io_in_bits_tc0_ot1_tg0_matrix_b),
    .io_in_bits_tc0_ot1_tg0_matrix_c(top_io_in_bits_tc0_ot1_tg0_matrix_c),
    .io_in_bits_tc0_ot1_tg4_matrix_a(top_io_in_bits_tc0_ot1_tg4_matrix_a),
    .io_in_bits_tc0_ot1_tg4_matrix_b(top_io_in_bits_tc0_ot1_tg4_matrix_b),
    .io_in_bits_tc0_ot1_tg4_matrix_c(top_io_in_bits_tc0_ot1_tg4_matrix_c),
    .io_in_bits_tc1_ot0_tg0_matrix_a(top_io_in_bits_tc1_ot0_tg0_matrix_a),
    .io_in_bits_tc1_ot0_tg0_matrix_b(top_io_in_bits_tc1_ot0_tg0_matrix_b),
    .io_in_bits_tc1_ot0_tg0_matrix_c(top_io_in_bits_tc1_ot0_tg0_matrix_c),
    .io_in_bits_tc1_ot0_tg4_matrix_a(top_io_in_bits_tc1_ot0_tg4_matrix_a),
    .io_in_bits_tc1_ot0_tg4_matrix_b(top_io_in_bits_tc1_ot0_tg4_matrix_b),
    .io_in_bits_tc1_ot0_tg4_matrix_c(top_io_in_bits_tc1_ot0_tg4_matrix_c),
    .io_in_bits_tc1_ot1_tg0_matrix_a(top_io_in_bits_tc1_ot1_tg0_matrix_a),
    .io_in_bits_tc1_ot1_tg0_matrix_b(top_io_in_bits_tc1_ot1_tg0_matrix_b),
    .io_in_bits_tc1_ot1_tg0_matrix_c(top_io_in_bits_tc1_ot1_tg0_matrix_c),
    .io_in_bits_tc1_ot1_tg4_matrix_a(top_io_in_bits_tc1_ot1_tg4_matrix_a),
    .io_in_bits_tc1_ot1_tg4_matrix_b(top_io_in_bits_tc1_ot1_tg4_matrix_b),
    .io_in_bits_tc1_ot1_tg4_matrix_c(top_io_in_bits_tc1_ot1_tg4_matrix_c),
    .io_in_bits_ctrl_matBSel(top_io_in_bits_ctrl_matBSel),
    .io_in_bits_ctrl_mixPcMode(top_io_in_bits_ctrl_mixPcMode),
    .io_out_valid(top_io_out_valid),
    .io_out_bits_tc0_octet0_threadgroup0_matrix_d_data(top_io_out_bits_tc0_octet0_threadgroup0_matrix_d_data),
    .io_out_bits_tc0_octet0_threadgroup4_matrix_d_data(top_io_out_bits_tc0_octet0_threadgroup4_matrix_d_data),
    .io_out_bits_tc0_octet1_threadgroup0_matrix_d_data(top_io_out_bits_tc0_octet1_threadgroup0_matrix_d_data),
    .io_out_bits_tc0_octet1_threadgroup4_matrix_d_data(top_io_out_bits_tc0_octet1_threadgroup4_matrix_d_data),
    .io_out_bits_tc1_octet0_threadgroup0_matrix_d_data(top_io_out_bits_tc1_octet0_threadgroup0_matrix_d_data),
    .io_out_bits_tc1_octet0_threadgroup4_matrix_d_data(top_io_out_bits_tc1_octet0_threadgroup4_matrix_d_data),
    .io_out_bits_tc1_octet1_threadgroup0_matrix_d_data(top_io_out_bits_tc1_octet1_threadgroup0_matrix_d_data),
    .io_out_bits_tc1_octet1_threadgroup4_matrix_d_data(top_io_out_bits_tc1_octet1_threadgroup4_matrix_d_data)
  );
  assign io_uart_ctrl_tx_en = manager_io_uart_ctrl_tx_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Adagio.scala 21:24]
  assign io_rf_r_data = manager_io_uart_rf_r_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Adagio.scala 25:22]
  assign manager_clock = clock;
  assign manager_reset = reset;
  assign manager_io_mixPc = io_mixPc; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Adagio.scala 27:20]
  assign manager_io_uart_ctrl_tx_done = io_uart_ctrl_tx_done; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Adagio.scala 21:24]
  assign manager_io_uart_ctrl_rx_valid = io_uart_ctrl_rx_valid; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Adagio.scala 21:24]
  assign manager_io_uart_rf_w_en = io_rf_w_en; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Adagio.scala 25:22]
  assign manager_io_uart_rf_r_addr = io_rf_r_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Adagio.scala 25:22]
  assign manager_io_uart_rf_w_addr = io_rf_w_addr; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Adagio.scala 25:22]
  assign manager_io_uart_rf_w_data = io_rf_w_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Adagio.scala 25:22]
  assign manager_io_top_src_ready = top_io_in_ready; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Adagio.scala 18:13]
  assign manager_io_top_wb_valid = top_io_out_valid; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Adagio.scala 19:21]
  assign manager_io_top_wb_bits_tc0_octet0_threadgroup0_matrix_d_data =
    top_io_out_bits_tc0_octet0_threadgroup0_matrix_d_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Adagio.scala 19:21]
  assign manager_io_top_wb_bits_tc0_octet0_threadgroup4_matrix_d_data =
    top_io_out_bits_tc0_octet0_threadgroup4_matrix_d_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Adagio.scala 19:21]
  assign manager_io_top_wb_bits_tc0_octet1_threadgroup0_matrix_d_data =
    top_io_out_bits_tc0_octet1_threadgroup0_matrix_d_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Adagio.scala 19:21]
  assign manager_io_top_wb_bits_tc0_octet1_threadgroup4_matrix_d_data =
    top_io_out_bits_tc0_octet1_threadgroup4_matrix_d_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Adagio.scala 19:21]
  assign manager_io_top_wb_bits_tc1_octet0_threadgroup0_matrix_d_data =
    top_io_out_bits_tc1_octet0_threadgroup0_matrix_d_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Adagio.scala 19:21]
  assign manager_io_top_wb_bits_tc1_octet0_threadgroup4_matrix_d_data =
    top_io_out_bits_tc1_octet0_threadgroup4_matrix_d_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Adagio.scala 19:21]
  assign manager_io_top_wb_bits_tc1_octet1_threadgroup0_matrix_d_data =
    top_io_out_bits_tc1_octet1_threadgroup0_matrix_d_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Adagio.scala 19:21]
  assign manager_io_top_wb_bits_tc1_octet1_threadgroup4_matrix_d_data =
    top_io_out_bits_tc1_octet1_threadgroup4_matrix_d_data; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Adagio.scala 19:21]
  assign top_clock = clock;
  assign top_reset = reset;
  assign top_io_in_valid = manager_io_top_src_valid; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Adagio.scala 18:13]
  assign top_io_in_bits_tc0_ot0_tg0_matrix_a = manager_io_top_src_bits_tc0_ot0_tg0_matrix_a; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Adagio.scala 18:13]
  assign top_io_in_bits_tc0_ot0_tg0_matrix_b = manager_io_top_src_bits_tc0_ot0_tg0_matrix_b; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Adagio.scala 18:13]
  assign top_io_in_bits_tc0_ot0_tg0_matrix_c = manager_io_top_src_bits_tc0_ot0_tg0_matrix_c; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Adagio.scala 18:13]
  assign top_io_in_bits_tc0_ot0_tg4_matrix_a = manager_io_top_src_bits_tc0_ot0_tg4_matrix_a; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Adagio.scala 18:13]
  assign top_io_in_bits_tc0_ot0_tg4_matrix_b = manager_io_top_src_bits_tc0_ot0_tg4_matrix_b; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Adagio.scala 18:13]
  assign top_io_in_bits_tc0_ot0_tg4_matrix_c = manager_io_top_src_bits_tc0_ot0_tg4_matrix_c; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Adagio.scala 18:13]
  assign top_io_in_bits_tc0_ot1_tg0_matrix_a = manager_io_top_src_bits_tc0_ot1_tg0_matrix_a; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Adagio.scala 18:13]
  assign top_io_in_bits_tc0_ot1_tg0_matrix_b = manager_io_top_src_bits_tc0_ot1_tg0_matrix_b; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Adagio.scala 18:13]
  assign top_io_in_bits_tc0_ot1_tg0_matrix_c = manager_io_top_src_bits_tc0_ot1_tg0_matrix_c; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Adagio.scala 18:13]
  assign top_io_in_bits_tc0_ot1_tg4_matrix_a = manager_io_top_src_bits_tc0_ot1_tg4_matrix_a; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Adagio.scala 18:13]
  assign top_io_in_bits_tc0_ot1_tg4_matrix_b = manager_io_top_src_bits_tc0_ot1_tg4_matrix_b; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Adagio.scala 18:13]
  assign top_io_in_bits_tc0_ot1_tg4_matrix_c = manager_io_top_src_bits_tc0_ot1_tg4_matrix_c; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Adagio.scala 18:13]
  assign top_io_in_bits_tc1_ot0_tg0_matrix_a = manager_io_top_src_bits_tc1_ot0_tg0_matrix_a; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Adagio.scala 18:13]
  assign top_io_in_bits_tc1_ot0_tg0_matrix_b = manager_io_top_src_bits_tc1_ot0_tg0_matrix_b; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Adagio.scala 18:13]
  assign top_io_in_bits_tc1_ot0_tg0_matrix_c = manager_io_top_src_bits_tc1_ot0_tg0_matrix_c; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Adagio.scala 18:13]
  assign top_io_in_bits_tc1_ot0_tg4_matrix_a = manager_io_top_src_bits_tc1_ot0_tg4_matrix_a; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Adagio.scala 18:13]
  assign top_io_in_bits_tc1_ot0_tg4_matrix_b = manager_io_top_src_bits_tc1_ot0_tg4_matrix_b; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Adagio.scala 18:13]
  assign top_io_in_bits_tc1_ot0_tg4_matrix_c = manager_io_top_src_bits_tc1_ot0_tg4_matrix_c; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Adagio.scala 18:13]
  assign top_io_in_bits_tc1_ot1_tg0_matrix_a = manager_io_top_src_bits_tc1_ot1_tg0_matrix_a; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Adagio.scala 18:13]
  assign top_io_in_bits_tc1_ot1_tg0_matrix_b = manager_io_top_src_bits_tc1_ot1_tg0_matrix_b; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Adagio.scala 18:13]
  assign top_io_in_bits_tc1_ot1_tg0_matrix_c = manager_io_top_src_bits_tc1_ot1_tg0_matrix_c; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Adagio.scala 18:13]
  assign top_io_in_bits_tc1_ot1_tg4_matrix_a = manager_io_top_src_bits_tc1_ot1_tg4_matrix_a; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Adagio.scala 18:13]
  assign top_io_in_bits_tc1_ot1_tg4_matrix_b = manager_io_top_src_bits_tc1_ot1_tg4_matrix_b; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Adagio.scala 18:13]
  assign top_io_in_bits_tc1_ot1_tg4_matrix_c = manager_io_top_src_bits_tc1_ot1_tg4_matrix_c; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Adagio.scala 18:13]
  assign top_io_in_bits_ctrl_matBSel = manager_io_top_src_bits_ctrl_matBSel; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Adagio.scala 18:13]
  assign top_io_in_bits_ctrl_mixPcMode = manager_io_top_src_bits_ctrl_mixPcMode; // @[Users/liuyuxuan/proc/Adagio/src/main/scala/System/Adagio.scala 18:13]
endmodule
